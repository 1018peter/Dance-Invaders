`include "constants.svh"
module level_pixel(
    input clk,
    input [LEVEL_SIZE-1:0] level,
    input [9:0] h_cnt,
    input [9:0] v_cnt,
    output logic [11:0] pixel_out,
    output logic valid
    );
    logic [5:0] mem_txt_addr;
    reg reg_h_cnt_compressed;
    reg reg_v_cnt_compressed;
parameter L=21;
parameter E=14;
parameter V=31;

always@* begin
    valid=0;
    mem_txt_addr=0;
    reg_h_cnt_compressed=0;
    reg_v_cnt_compressed=0;
    if(v_cnt>=28&&v_cnt<140) begin
            if(h_cnt>=120&&h_cnt<200) begin
            mem_txt_addr=L;
            reg_h_cnt_compressed=(h_cnt-120)>>4;
            reg_v_cnt_compressed=(v_cnt-28)>>4;
            valid=1;
            end
            else if(h_cnt>=200&&h_cnt<280) begin
            reg_h_cnt_compressed=(h_cnt-200)>>4;
            reg_v_cnt_compressed=(v_cnt-28)>>4;
            mem_txt_addr=E;
            valid=1;
            end
            else if(h_cnt>=280&&h_cnt<360) begin
            mem_txt_addr=V;
            reg_h_cnt_compressed=(h_cnt-280)>>4;
            reg_v_cnt_compressed=(v_cnt-28)>>4;
            valid=1;
            end
            else if(h_cnt>=360&&h_cnt<440)begin
            mem_txt_addr=E;
            reg_h_cnt_compressed=(h_cnt-360)>>4;
            reg_v_cnt_compressed=(v_cnt-28)>>4;
            valid=1;
            end
            else if(h_cnt>=440&&h_cnt<520)begin
            mem_txt_addr=L;
            reg_h_cnt_compressed=(h_cnt-440)>>4;
            reg_v_cnt_compressed=(v_cnt-28)>>4;
            valid=1;
            end
        end

        else if(v_cnt>=160&&v_cnt<272) begin
            if(h_cnt>=240&&h_cnt<320) begin
            reg_h_cnt_compressed=(h_cnt-240)>>4;
            reg_v_cnt_compressed=(v_cnt-160)>>4;
            mem_txt_addr=level/10;
            valid=1;
        end
        else if(h_cnt>=320&&h_cnt<400) begin
            mem_txt_addr=level%10;
            reg_h_cnt_compressed=(h_cnt-320)>>4;
            reg_v_cnt_compressed=(v_cnt-160)>>4;
            valid=1;
        end

        end
end
        memory_txt level_show(
        .clk(clk),
        .txt_addr(mem_txt_addr),
        .h_point(wire_h_cnt_compressed),
        .v_point(wire_v_cnt_compressed),
        .pixel(pixel_out)
    );

endmodule

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/01/02 13:57:31
// Design Name: 
// Module Name: alien_pixel_reader
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module alien_pixel_reader(
    input [1:0] frame_num,
    input [1:0] alien_type,
    input [3:0] size_select,
    input [1:0] deriv_select,
    input [15:0] pixel_addr,
    output logic palette_out
    );
    
    
reg size0_type0_frame0_deriv0 [0:2047];
reg size0_type0_frame0_deriv1 [0:2047];
reg size0_type0_frame0_deriv2 [0:2047];
reg size0_type0_frame0_deriv3 [0:2047];
reg size0_type0_frame1_deriv0 [0:2047];
reg size0_type0_frame1_deriv1 [0:2047];
reg size0_type0_frame1_deriv2 [0:2047];
reg size0_type0_frame1_deriv3 [0:2047];
reg size0_type1_frame0_deriv0 [0:2047];
reg size0_type1_frame0_deriv1 [0:2047];
reg size0_type1_frame0_deriv2 [0:2047];
reg size0_type1_frame0_deriv3 [0:2047];
reg size0_type1_frame1_deriv0 [0:2047];
reg size0_type1_frame1_deriv1 [0:2047];
reg size0_type1_frame1_deriv2 [0:2047];
reg size0_type1_frame1_deriv3 [0:2047];
reg size1_type0_frame0_deriv0 [0:1921];
reg size1_type0_frame0_deriv1 [0:1921];
reg size1_type0_frame0_deriv2 [0:1921];
reg size1_type0_frame0_deriv3 [0:1921];
reg size1_type0_frame1_deriv0 [0:1921];
reg size1_type0_frame1_deriv1 [0:1921];
reg size1_type0_frame1_deriv2 [0:1921];
reg size1_type0_frame1_deriv3 [0:1921];
reg size1_type1_frame0_deriv0 [0:1921];
reg size1_type1_frame0_deriv1 [0:1921];
reg size1_type1_frame0_deriv2 [0:1921];
reg size1_type1_frame0_deriv3 [0:1921];
reg size1_type1_frame1_deriv0 [0:1921];
reg size1_type1_frame1_deriv1 [0:1921];
reg size1_type1_frame1_deriv2 [0:1921];
reg size1_type1_frame1_deriv3 [0:1921];
reg size2_type0_frame0_deriv0 [0:1799];
reg size2_type0_frame0_deriv1 [0:1799];
reg size2_type0_frame0_deriv2 [0:1799];
reg size2_type0_frame0_deriv3 [0:1799];
reg size2_type0_frame1_deriv0 [0:1799];
reg size2_type0_frame1_deriv1 [0:1799];
reg size2_type0_frame1_deriv2 [0:1799];
reg size2_type0_frame1_deriv3 [0:1799];
reg size2_type1_frame0_deriv0 [0:1799];
reg size2_type1_frame0_deriv1 [0:1799];
reg size2_type1_frame0_deriv2 [0:1799];
reg size2_type1_frame0_deriv3 [0:1799];
reg size2_type1_frame1_deriv0 [0:1799];
reg size2_type1_frame1_deriv1 [0:1799];
reg size2_type1_frame1_deriv2 [0:1799];
reg size2_type1_frame1_deriv3 [0:1799];
reg size3_type0_frame0_deriv0 [0:1681];
reg size3_type0_frame0_deriv1 [0:1681];
reg size3_type0_frame0_deriv2 [0:1681];
reg size3_type0_frame0_deriv3 [0:1681];
reg size3_type0_frame1_deriv0 [0:1681];
reg size3_type0_frame1_deriv1 [0:1681];
reg size3_type0_frame1_deriv2 [0:1681];
reg size3_type0_frame1_deriv3 [0:1681];
reg size3_type1_frame0_deriv0 [0:1681];
reg size3_type1_frame0_deriv1 [0:1681];
reg size3_type1_frame0_deriv2 [0:1681];
reg size3_type1_frame0_deriv3 [0:1681];
reg size3_type1_frame1_deriv0 [0:1681];
reg size3_type1_frame1_deriv1 [0:1681];
reg size3_type1_frame1_deriv2 [0:1681];
reg size3_type1_frame1_deriv3 [0:1681];
reg size4_type0_frame0_deriv0 [0:1567];
reg size4_type0_frame0_deriv1 [0:1567];
reg size4_type0_frame0_deriv2 [0:1567];
reg size4_type0_frame0_deriv3 [0:1567];
reg size4_type0_frame1_deriv0 [0:1567];
reg size4_type0_frame1_deriv1 [0:1567];
reg size4_type0_frame1_deriv2 [0:1567];
reg size4_type0_frame1_deriv3 [0:1567];
reg size4_type1_frame0_deriv0 [0:1567];
reg size4_type1_frame0_deriv1 [0:1567];
reg size4_type1_frame0_deriv2 [0:1567];
reg size4_type1_frame0_deriv3 [0:1567];
reg size4_type1_frame1_deriv0 [0:1567];
reg size4_type1_frame1_deriv1 [0:1567];
reg size4_type1_frame1_deriv2 [0:1567];
reg size4_type1_frame1_deriv3 [0:1567];
reg size5_type0_frame0_deriv0 [0:1457];
reg size5_type0_frame0_deriv1 [0:1457];
reg size5_type0_frame0_deriv2 [0:1457];
reg size5_type0_frame0_deriv3 [0:1457];
reg size5_type0_frame1_deriv0 [0:1457];
reg size5_type0_frame1_deriv1 [0:1457];
reg size5_type0_frame1_deriv2 [0:1457];
reg size5_type0_frame1_deriv3 [0:1457];
reg size5_type1_frame0_deriv0 [0:1457];
reg size5_type1_frame0_deriv1 [0:1457];
reg size5_type1_frame0_deriv2 [0:1457];
reg size5_type1_frame0_deriv3 [0:1457];
reg size5_type1_frame1_deriv0 [0:1457];
reg size5_type1_frame1_deriv1 [0:1457];
reg size5_type1_frame1_deriv2 [0:1457];
reg size5_type1_frame1_deriv3 [0:1457];
reg size6_type0_frame0_deriv0 [0:1351];
reg size6_type0_frame0_deriv1 [0:1351];
reg size6_type0_frame0_deriv2 [0:1351];
reg size6_type0_frame0_deriv3 [0:1351];
reg size6_type0_frame1_deriv0 [0:1351];
reg size6_type0_frame1_deriv1 [0:1351];
reg size6_type0_frame1_deriv2 [0:1351];
reg size6_type0_frame1_deriv3 [0:1351];
reg size6_type1_frame0_deriv0 [0:1351];
reg size6_type1_frame0_deriv1 [0:1351];
reg size6_type1_frame0_deriv2 [0:1351];
reg size6_type1_frame0_deriv3 [0:1351];
reg size6_type1_frame1_deriv0 [0:1351];
reg size6_type1_frame1_deriv1 [0:1351];
reg size6_type1_frame1_deriv2 [0:1351];
reg size6_type1_frame1_deriv3 [0:1351];
reg size7_type0_frame0_deriv0 [0:1249];
reg size7_type0_frame0_deriv1 [0:1249];
reg size7_type0_frame0_deriv2 [0:1249];
reg size7_type0_frame0_deriv3 [0:1249];
reg size7_type0_frame1_deriv0 [0:1249];
reg size7_type0_frame1_deriv1 [0:1249];
reg size7_type0_frame1_deriv2 [0:1249];
reg size7_type0_frame1_deriv3 [0:1249];
reg size7_type1_frame0_deriv0 [0:1249];
reg size7_type1_frame0_deriv1 [0:1249];
reg size7_type1_frame0_deriv2 [0:1249];
reg size7_type1_frame0_deriv3 [0:1249];
reg size7_type1_frame1_deriv0 [0:1249];
reg size7_type1_frame1_deriv1 [0:1249];
reg size7_type1_frame1_deriv2 [0:1249];
reg size7_type1_frame1_deriv3 [0:1249];
reg size8_type0_frame0_deriv0 [0:1151];
reg size8_type0_frame0_deriv1 [0:1151];
reg size8_type0_frame0_deriv2 [0:1151];
reg size8_type0_frame0_deriv3 [0:1151];
reg size8_type0_frame1_deriv0 [0:1151];
reg size8_type0_frame1_deriv1 [0:1151];
reg size8_type0_frame1_deriv2 [0:1151];
reg size8_type0_frame1_deriv3 [0:1151];
reg size8_type1_frame0_deriv0 [0:1151];
reg size8_type1_frame0_deriv1 [0:1151];
reg size8_type1_frame0_deriv2 [0:1151];
reg size8_type1_frame0_deriv3 [0:1151];
reg size8_type1_frame1_deriv0 [0:1151];
reg size8_type1_frame1_deriv1 [0:1151];
reg size8_type1_frame1_deriv2 [0:1151];
reg size8_type1_frame1_deriv3 [0:1151];
reg size9_type0_frame0_deriv0 [0:1057];
reg size9_type0_frame0_deriv1 [0:1057];
reg size9_type0_frame0_deriv2 [0:1057];
reg size9_type0_frame0_deriv3 [0:1057];
reg size9_type0_frame1_deriv0 [0:1057];
reg size9_type0_frame1_deriv1 [0:1057];
reg size9_type0_frame1_deriv2 [0:1057];
reg size9_type0_frame1_deriv3 [0:1057];
reg size9_type1_frame0_deriv0 [0:1057];
reg size9_type1_frame0_deriv1 [0:1057];
reg size9_type1_frame0_deriv2 [0:1057];
reg size9_type1_frame0_deriv3 [0:1057];
reg size9_type1_frame1_deriv0 [0:1057];
reg size9_type1_frame1_deriv1 [0:1057];
reg size9_type1_frame1_deriv2 [0:1057];
reg size9_type1_frame1_deriv3 [0:1057];
reg size10_type0_frame0_deriv0 [0:967];
reg size10_type0_frame0_deriv1 [0:967];
reg size10_type0_frame0_deriv2 [0:967];
reg size10_type0_frame0_deriv3 [0:967];
reg size10_type0_frame1_deriv0 [0:967];
reg size10_type0_frame1_deriv1 [0:967];
reg size10_type0_frame1_deriv2 [0:967];
reg size10_type0_frame1_deriv3 [0:967];
reg size10_type1_frame0_deriv0 [0:967];
reg size10_type1_frame0_deriv1 [0:967];
reg size10_type1_frame0_deriv2 [0:967];
reg size10_type1_frame0_deriv3 [0:967];
reg size10_type1_frame1_deriv0 [0:967];
reg size10_type1_frame1_deriv1 [0:967];
reg size10_type1_frame1_deriv2 [0:967];
reg size10_type1_frame1_deriv3 [0:967];
reg size11_type0_frame0_deriv0 [0:881];
reg size11_type0_frame0_deriv1 [0:881];
reg size11_type0_frame0_deriv2 [0:881];
reg size11_type0_frame0_deriv3 [0:881];
reg size11_type0_frame1_deriv0 [0:881];
reg size11_type0_frame1_deriv1 [0:881];
reg size11_type0_frame1_deriv2 [0:881];
reg size11_type0_frame1_deriv3 [0:881];
reg size11_type1_frame0_deriv0 [0:881];
reg size11_type1_frame0_deriv1 [0:881];
reg size11_type1_frame0_deriv2 [0:881];
reg size11_type1_frame0_deriv3 [0:881];
reg size11_type1_frame1_deriv0 [0:881];
reg size11_type1_frame1_deriv1 [0:881];
reg size11_type1_frame1_deriv2 [0:881];
reg size11_type1_frame1_deriv3 [0:881];
reg size12_type0_frame0_deriv0 [0:799];
reg size12_type0_frame0_deriv1 [0:799];
reg size12_type0_frame0_deriv2 [0:799];
reg size12_type0_frame0_deriv3 [0:799];
reg size12_type0_frame1_deriv0 [0:799];
reg size12_type0_frame1_deriv1 [0:799];
reg size12_type0_frame1_deriv2 [0:799];
reg size12_type0_frame1_deriv3 [0:799];
reg size12_type1_frame0_deriv0 [0:799];
reg size12_type1_frame0_deriv1 [0:799];
reg size12_type1_frame0_deriv2 [0:799];
reg size12_type1_frame0_deriv3 [0:799];
reg size12_type1_frame1_deriv0 [0:799];
reg size12_type1_frame1_deriv1 [0:799];
reg size12_type1_frame1_deriv2 [0:799];
reg size12_type1_frame1_deriv3 [0:799];
reg size13_type0_frame0_deriv0 [0:721];
reg size13_type0_frame0_deriv1 [0:721];
reg size13_type0_frame0_deriv2 [0:721];
reg size13_type0_frame0_deriv3 [0:721];
reg size13_type0_frame1_deriv0 [0:721];
reg size13_type0_frame1_deriv1 [0:721];
reg size13_type0_frame1_deriv2 [0:721];
reg size13_type0_frame1_deriv3 [0:721];
reg size13_type1_frame0_deriv0 [0:721];
reg size13_type1_frame0_deriv1 [0:721];
reg size13_type1_frame0_deriv2 [0:721];
reg size13_type1_frame0_deriv3 [0:721];
reg size13_type1_frame1_deriv0 [0:721];
reg size13_type1_frame1_deriv1 [0:721];
reg size13_type1_frame1_deriv2 [0:721];
reg size13_type1_frame1_deriv3 [0:721];
reg size14_type0_frame0_deriv0 [0:647];
reg size14_type0_frame0_deriv1 [0:647];
reg size14_type0_frame0_deriv2 [0:647];
reg size14_type0_frame0_deriv3 [0:647];
reg size14_type0_frame1_deriv0 [0:647];
reg size14_type0_frame1_deriv1 [0:647];
reg size14_type0_frame1_deriv2 [0:647];
reg size14_type0_frame1_deriv3 [0:647];
reg size14_type1_frame0_deriv0 [0:647];
reg size14_type1_frame0_deriv1 [0:647];
reg size14_type1_frame0_deriv2 [0:647];
reg size14_type1_frame0_deriv3 [0:647];
reg size14_type1_frame1_deriv0 [0:647];
reg size14_type1_frame1_deriv1 [0:647];
reg size14_type1_frame1_deriv2 [0:647];
reg size14_type1_frame1_deriv3 [0:647];
reg size15_type0_frame0_deriv0 [0:577];
reg size15_type0_frame0_deriv1 [0:577];
reg size15_type0_frame0_deriv2 [0:577];
reg size15_type0_frame0_deriv3 [0:577];
reg size15_type0_frame1_deriv0 [0:577];
reg size15_type0_frame1_deriv1 [0:577];
reg size15_type0_frame1_deriv2 [0:577];
reg size15_type0_frame1_deriv3 [0:577];
reg size15_type1_frame0_deriv0 [0:577];
reg size15_type1_frame0_deriv1 [0:577];
reg size15_type1_frame0_deriv2 [0:577];
reg size15_type1_frame0_deriv3 [0:577];
reg size15_type1_frame1_deriv0 [0:577];
reg size15_type1_frame1_deriv1 [0:577];
reg size15_type1_frame1_deriv2 [0:577];
reg size15_type1_frame1_deriv3 [0:577];


initial begin
$readmemb("size0_type0_frame0_deriv0.mem", size0_type0_frame0_deriv0);
$readmemb("size0_type0_frame0_deriv1.mem", size0_type0_frame0_deriv1);
$readmemb("size0_type0_frame0_deriv2.mem", size0_type0_frame0_deriv2);
$readmemb("size0_type0_frame0_deriv3.mem", size0_type0_frame0_deriv3);
$readmemb("size0_type0_frame1_deriv0.mem", size0_type0_frame1_deriv0);
$readmemb("size0_type0_frame1_deriv1.mem", size0_type0_frame1_deriv1);
$readmemb("size0_type0_frame1_deriv2.mem", size0_type0_frame1_deriv2);
$readmemb("size0_type0_frame1_deriv3.mem", size0_type0_frame1_deriv3);
$readmemb("size0_type1_frame0_deriv0.mem", size0_type1_frame0_deriv0);
$readmemb("size0_type1_frame0_deriv1.mem", size0_type1_frame0_deriv1);
$readmemb("size0_type1_frame0_deriv2.mem", size0_type1_frame0_deriv2);
$readmemb("size0_type1_frame0_deriv3.mem", size0_type1_frame0_deriv3);
$readmemb("size0_type1_frame1_deriv0.mem", size0_type1_frame1_deriv0);
$readmemb("size0_type1_frame1_deriv1.mem", size0_type1_frame1_deriv1);
$readmemb("size0_type1_frame1_deriv2.mem", size0_type1_frame1_deriv2);
$readmemb("size0_type1_frame1_deriv3.mem", size0_type1_frame1_deriv3);
$readmemb("size1_type0_frame0_deriv0.mem", size1_type0_frame0_deriv0);
$readmemb("size1_type0_frame0_deriv1.mem", size1_type0_frame0_deriv1);
$readmemb("size1_type0_frame0_deriv2.mem", size1_type0_frame0_deriv2);
$readmemb("size1_type0_frame0_deriv3.mem", size1_type0_frame0_deriv3);
$readmemb("size1_type0_frame1_deriv0.mem", size1_type0_frame1_deriv0);
$readmemb("size1_type0_frame1_deriv1.mem", size1_type0_frame1_deriv1);
$readmemb("size1_type0_frame1_deriv2.mem", size1_type0_frame1_deriv2);
$readmemb("size1_type0_frame1_deriv3.mem", size1_type0_frame1_deriv3);
$readmemb("size1_type1_frame0_deriv0.mem", size1_type1_frame0_deriv0);
$readmemb("size1_type1_frame0_deriv1.mem", size1_type1_frame0_deriv1);
$readmemb("size1_type1_frame0_deriv2.mem", size1_type1_frame0_deriv2);
$readmemb("size1_type1_frame0_deriv3.mem", size1_type1_frame0_deriv3);
$readmemb("size1_type1_frame1_deriv0.mem", size1_type1_frame1_deriv0);
$readmemb("size1_type1_frame1_deriv1.mem", size1_type1_frame1_deriv1);
$readmemb("size1_type1_frame1_deriv2.mem", size1_type1_frame1_deriv2);
$readmemb("size1_type1_frame1_deriv3.mem", size1_type1_frame1_deriv3);
$readmemb("size2_type0_frame0_deriv0.mem", size2_type0_frame0_deriv0);
$readmemb("size2_type0_frame0_deriv1.mem", size2_type0_frame0_deriv1);
$readmemb("size2_type0_frame0_deriv2.mem", size2_type0_frame0_deriv2);
$readmemb("size2_type0_frame0_deriv3.mem", size2_type0_frame0_deriv3);
$readmemb("size2_type0_frame1_deriv0.mem", size2_type0_frame1_deriv0);
$readmemb("size2_type0_frame1_deriv1.mem", size2_type0_frame1_deriv1);
$readmemb("size2_type0_frame1_deriv2.mem", size2_type0_frame1_deriv2);
$readmemb("size2_type0_frame1_deriv3.mem", size2_type0_frame1_deriv3);
$readmemb("size2_type1_frame0_deriv0.mem", size2_type1_frame0_deriv0);
$readmemb("size2_type1_frame0_deriv1.mem", size2_type1_frame0_deriv1);
$readmemb("size2_type1_frame0_deriv2.mem", size2_type1_frame0_deriv2);
$readmemb("size2_type1_frame0_deriv3.mem", size2_type1_frame0_deriv3);
$readmemb("size2_type1_frame1_deriv0.mem", size2_type1_frame1_deriv0);
$readmemb("size2_type1_frame1_deriv1.mem", size2_type1_frame1_deriv1);
$readmemb("size2_type1_frame1_deriv2.mem", size2_type1_frame1_deriv2);
$readmemb("size2_type1_frame1_deriv3.mem", size2_type1_frame1_deriv3);
$readmemb("size3_type0_frame0_deriv0.mem", size3_type0_frame0_deriv0);
$readmemb("size3_type0_frame0_deriv1.mem", size3_type0_frame0_deriv1);
$readmemb("size3_type0_frame0_deriv2.mem", size3_type0_frame0_deriv2);
$readmemb("size3_type0_frame0_deriv3.mem", size3_type0_frame0_deriv3);
$readmemb("size3_type0_frame1_deriv0.mem", size3_type0_frame1_deriv0);
$readmemb("size3_type0_frame1_deriv1.mem", size3_type0_frame1_deriv1);
$readmemb("size3_type0_frame1_deriv2.mem", size3_type0_frame1_deriv2);
$readmemb("size3_type0_frame1_deriv3.mem", size3_type0_frame1_deriv3);
$readmemb("size3_type1_frame0_deriv0.mem", size3_type1_frame0_deriv0);
$readmemb("size3_type1_frame0_deriv1.mem", size3_type1_frame0_deriv1);
$readmemb("size3_type1_frame0_deriv2.mem", size3_type1_frame0_deriv2);
$readmemb("size3_type1_frame0_deriv3.mem", size3_type1_frame0_deriv3);
$readmemb("size3_type1_frame1_deriv0.mem", size3_type1_frame1_deriv0);
$readmemb("size3_type1_frame1_deriv1.mem", size3_type1_frame1_deriv1);
$readmemb("size3_type1_frame1_deriv2.mem", size3_type1_frame1_deriv2);
$readmemb("size3_type1_frame1_deriv3.mem", size3_type1_frame1_deriv3);
$readmemb("size4_type0_frame0_deriv0.mem", size4_type0_frame0_deriv0);
$readmemb("size4_type0_frame0_deriv1.mem", size4_type0_frame0_deriv1);
$readmemb("size4_type0_frame0_deriv2.mem", size4_type0_frame0_deriv2);
$readmemb("size4_type0_frame0_deriv3.mem", size4_type0_frame0_deriv3);
$readmemb("size4_type0_frame1_deriv0.mem", size4_type0_frame1_deriv0);
$readmemb("size4_type0_frame1_deriv1.mem", size4_type0_frame1_deriv1);
$readmemb("size4_type0_frame1_deriv2.mem", size4_type0_frame1_deriv2);
$readmemb("size4_type0_frame1_deriv3.mem", size4_type0_frame1_deriv3);
$readmemb("size4_type1_frame0_deriv0.mem", size4_type1_frame0_deriv0);
$readmemb("size4_type1_frame0_deriv1.mem", size4_type1_frame0_deriv1);
$readmemb("size4_type1_frame0_deriv2.mem", size4_type1_frame0_deriv2);
$readmemb("size4_type1_frame0_deriv3.mem", size4_type1_frame0_deriv3);
$readmemb("size4_type1_frame1_deriv0.mem", size4_type1_frame1_deriv0);
$readmemb("size4_type1_frame1_deriv1.mem", size4_type1_frame1_deriv1);
$readmemb("size4_type1_frame1_deriv2.mem", size4_type1_frame1_deriv2);
$readmemb("size4_type1_frame1_deriv3.mem", size4_type1_frame1_deriv3);
$readmemb("size5_type0_frame0_deriv0.mem", size5_type0_frame0_deriv0);
$readmemb("size5_type0_frame0_deriv1.mem", size5_type0_frame0_deriv1);
$readmemb("size5_type0_frame0_deriv2.mem", size5_type0_frame0_deriv2);
$readmemb("size5_type0_frame0_deriv3.mem", size5_type0_frame0_deriv3);
$readmemb("size5_type0_frame1_deriv0.mem", size5_type0_frame1_deriv0);
$readmemb("size5_type0_frame1_deriv1.mem", size5_type0_frame1_deriv1);
$readmemb("size5_type0_frame1_deriv2.mem", size5_type0_frame1_deriv2);
$readmemb("size5_type0_frame1_deriv3.mem", size5_type0_frame1_deriv3);
$readmemb("size5_type1_frame0_deriv0.mem", size5_type1_frame0_deriv0);
$readmemb("size5_type1_frame0_deriv1.mem", size5_type1_frame0_deriv1);
$readmemb("size5_type1_frame0_deriv2.mem", size5_type1_frame0_deriv2);
$readmemb("size5_type1_frame0_deriv3.mem", size5_type1_frame0_deriv3);
$readmemb("size5_type1_frame1_deriv0.mem", size5_type1_frame1_deriv0);
$readmemb("size5_type1_frame1_deriv1.mem", size5_type1_frame1_deriv1);
$readmemb("size5_type1_frame1_deriv2.mem", size5_type1_frame1_deriv2);
$readmemb("size5_type1_frame1_deriv3.mem", size5_type1_frame1_deriv3);
$readmemb("size6_type0_frame0_deriv0.mem", size6_type0_frame0_deriv0);
$readmemb("size6_type0_frame0_deriv1.mem", size6_type0_frame0_deriv1);
$readmemb("size6_type0_frame0_deriv2.mem", size6_type0_frame0_deriv2);
$readmemb("size6_type0_frame0_deriv3.mem", size6_type0_frame0_deriv3);
$readmemb("size6_type0_frame1_deriv0.mem", size6_type0_frame1_deriv0);
$readmemb("size6_type0_frame1_deriv1.mem", size6_type0_frame1_deriv1);
$readmemb("size6_type0_frame1_deriv2.mem", size6_type0_frame1_deriv2);
$readmemb("size6_type0_frame1_deriv3.mem", size6_type0_frame1_deriv3);
$readmemb("size6_type1_frame0_deriv0.mem", size6_type1_frame0_deriv0);
$readmemb("size6_type1_frame0_deriv1.mem", size6_type1_frame0_deriv1);
$readmemb("size6_type1_frame0_deriv2.mem", size6_type1_frame0_deriv2);
$readmemb("size6_type1_frame0_deriv3.mem", size6_type1_frame0_deriv3);
$readmemb("size6_type1_frame1_deriv0.mem", size6_type1_frame1_deriv0);
$readmemb("size6_type1_frame1_deriv1.mem", size6_type1_frame1_deriv1);
$readmemb("size6_type1_frame1_deriv2.mem", size6_type1_frame1_deriv2);
$readmemb("size6_type1_frame1_deriv3.mem", size6_type1_frame1_deriv3);
$readmemb("size7_type0_frame0_deriv0.mem", size7_type0_frame0_deriv0);
$readmemb("size7_type0_frame0_deriv1.mem", size7_type0_frame0_deriv1);
$readmemb("size7_type0_frame0_deriv2.mem", size7_type0_frame0_deriv2);
$readmemb("size7_type0_frame0_deriv3.mem", size7_type0_frame0_deriv3);
$readmemb("size7_type0_frame1_deriv0.mem", size7_type0_frame1_deriv0);
$readmemb("size7_type0_frame1_deriv1.mem", size7_type0_frame1_deriv1);
$readmemb("size7_type0_frame1_deriv2.mem", size7_type0_frame1_deriv2);
$readmemb("size7_type0_frame1_deriv3.mem", size7_type0_frame1_deriv3);
$readmemb("size7_type1_frame0_deriv0.mem", size7_type1_frame0_deriv0);
$readmemb("size7_type1_frame0_deriv1.mem", size7_type1_frame0_deriv1);
$readmemb("size7_type1_frame0_deriv2.mem", size7_type1_frame0_deriv2);
$readmemb("size7_type1_frame0_deriv3.mem", size7_type1_frame0_deriv3);
$readmemb("size7_type1_frame1_deriv0.mem", size7_type1_frame1_deriv0);
$readmemb("size7_type1_frame1_deriv1.mem", size7_type1_frame1_deriv1);
$readmemb("size7_type1_frame1_deriv2.mem", size7_type1_frame1_deriv2);
$readmemb("size7_type1_frame1_deriv3.mem", size7_type1_frame1_deriv3);
$readmemb("size8_type0_frame0_deriv0.mem", size8_type0_frame0_deriv0);
$readmemb("size8_type0_frame0_deriv1.mem", size8_type0_frame0_deriv1);
$readmemb("size8_type0_frame0_deriv2.mem", size8_type0_frame0_deriv2);
$readmemb("size8_type0_frame0_deriv3.mem", size8_type0_frame0_deriv3);
$readmemb("size8_type0_frame1_deriv0.mem", size8_type0_frame1_deriv0);
$readmemb("size8_type0_frame1_deriv1.mem", size8_type0_frame1_deriv1);
$readmemb("size8_type0_frame1_deriv2.mem", size8_type0_frame1_deriv2);
$readmemb("size8_type0_frame1_deriv3.mem", size8_type0_frame1_deriv3);
$readmemb("size8_type1_frame0_deriv0.mem", size8_type1_frame0_deriv0);
$readmemb("size8_type1_frame0_deriv1.mem", size8_type1_frame0_deriv1);
$readmemb("size8_type1_frame0_deriv2.mem", size8_type1_frame0_deriv2);
$readmemb("size8_type1_frame0_deriv3.mem", size8_type1_frame0_deriv3);
$readmemb("size8_type1_frame1_deriv0.mem", size8_type1_frame1_deriv0);
$readmemb("size8_type1_frame1_deriv1.mem", size8_type1_frame1_deriv1);
$readmemb("size8_type1_frame1_deriv2.mem", size8_type1_frame1_deriv2);
$readmemb("size8_type1_frame1_deriv3.mem", size8_type1_frame1_deriv3);
$readmemb("size9_type0_frame0_deriv0.mem", size9_type0_frame0_deriv0);
$readmemb("size9_type0_frame0_deriv1.mem", size9_type0_frame0_deriv1);
$readmemb("size9_type0_frame0_deriv2.mem", size9_type0_frame0_deriv2);
$readmemb("size9_type0_frame0_deriv3.mem", size9_type0_frame0_deriv3);
$readmemb("size9_type0_frame1_deriv0.mem", size9_type0_frame1_deriv0);
$readmemb("size9_type0_frame1_deriv1.mem", size9_type0_frame1_deriv1);
$readmemb("size9_type0_frame1_deriv2.mem", size9_type0_frame1_deriv2);
$readmemb("size9_type0_frame1_deriv3.mem", size9_type0_frame1_deriv3);
$readmemb("size9_type1_frame0_deriv0.mem", size9_type1_frame0_deriv0);
$readmemb("size9_type1_frame0_deriv1.mem", size9_type1_frame0_deriv1);
$readmemb("size9_type1_frame0_deriv2.mem", size9_type1_frame0_deriv2);
$readmemb("size9_type1_frame0_deriv3.mem", size9_type1_frame0_deriv3);
$readmemb("size9_type1_frame1_deriv0.mem", size9_type1_frame1_deriv0);
$readmemb("size9_type1_frame1_deriv1.mem", size9_type1_frame1_deriv1);
$readmemb("size9_type1_frame1_deriv2.mem", size9_type1_frame1_deriv2);
$readmemb("size9_type1_frame1_deriv3.mem", size9_type1_frame1_deriv3);
$readmemb("size10_type0_frame0_deriv0.mem", size10_type0_frame0_deriv0);
$readmemb("size10_type0_frame0_deriv1.mem", size10_type0_frame0_deriv1);
$readmemb("size10_type0_frame0_deriv2.mem", size10_type0_frame0_deriv2);
$readmemb("size10_type0_frame0_deriv3.mem", size10_type0_frame0_deriv3);
$readmemb("size10_type0_frame1_deriv0.mem", size10_type0_frame1_deriv0);
$readmemb("size10_type0_frame1_deriv1.mem", size10_type0_frame1_deriv1);
$readmemb("size10_type0_frame1_deriv2.mem", size10_type0_frame1_deriv2);
$readmemb("size10_type0_frame1_deriv3.mem", size10_type0_frame1_deriv3);
$readmemb("size10_type1_frame0_deriv0.mem", size10_type1_frame0_deriv0);
$readmemb("size10_type1_frame0_deriv1.mem", size10_type1_frame0_deriv1);
$readmemb("size10_type1_frame0_deriv2.mem", size10_type1_frame0_deriv2);
$readmemb("size10_type1_frame0_deriv3.mem", size10_type1_frame0_deriv3);
$readmemb("size10_type1_frame1_deriv0.mem", size10_type1_frame1_deriv0);
$readmemb("size10_type1_frame1_deriv1.mem", size10_type1_frame1_deriv1);
$readmemb("size10_type1_frame1_deriv2.mem", size10_type1_frame1_deriv2);
$readmemb("size10_type1_frame1_deriv3.mem", size10_type1_frame1_deriv3);
$readmemb("size11_type0_frame0_deriv0.mem", size11_type0_frame0_deriv0);
$readmemb("size11_type0_frame0_deriv1.mem", size11_type0_frame0_deriv1);
$readmemb("size11_type0_frame0_deriv2.mem", size11_type0_frame0_deriv2);
$readmemb("size11_type0_frame0_deriv3.mem", size11_type0_frame0_deriv3);
$readmemb("size11_type0_frame1_deriv0.mem", size11_type0_frame1_deriv0);
$readmemb("size11_type0_frame1_deriv1.mem", size11_type0_frame1_deriv1);
$readmemb("size11_type0_frame1_deriv2.mem", size11_type0_frame1_deriv2);
$readmemb("size11_type0_frame1_deriv3.mem", size11_type0_frame1_deriv3);
$readmemb("size11_type1_frame0_deriv0.mem", size11_type1_frame0_deriv0);
$readmemb("size11_type1_frame0_deriv1.mem", size11_type1_frame0_deriv1);
$readmemb("size11_type1_frame0_deriv2.mem", size11_type1_frame0_deriv2);
$readmemb("size11_type1_frame0_deriv3.mem", size11_type1_frame0_deriv3);
$readmemb("size11_type1_frame1_deriv0.mem", size11_type1_frame1_deriv0);
$readmemb("size11_type1_frame1_deriv1.mem", size11_type1_frame1_deriv1);
$readmemb("size11_type1_frame1_deriv2.mem", size11_type1_frame1_deriv2);
$readmemb("size11_type1_frame1_deriv3.mem", size11_type1_frame1_deriv3);
$readmemb("size12_type0_frame0_deriv0.mem", size12_type0_frame0_deriv0);
$readmemb("size12_type0_frame0_deriv1.mem", size12_type0_frame0_deriv1);
$readmemb("size12_type0_frame0_deriv2.mem", size12_type0_frame0_deriv2);
$readmemb("size12_type0_frame0_deriv3.mem", size12_type0_frame0_deriv3);
$readmemb("size12_type0_frame1_deriv0.mem", size12_type0_frame1_deriv0);
$readmemb("size12_type0_frame1_deriv1.mem", size12_type0_frame1_deriv1);
$readmemb("size12_type0_frame1_deriv2.mem", size12_type0_frame1_deriv2);
$readmemb("size12_type0_frame1_deriv3.mem", size12_type0_frame1_deriv3);
$readmemb("size12_type1_frame0_deriv0.mem", size12_type1_frame0_deriv0);
$readmemb("size12_type1_frame0_deriv1.mem", size12_type1_frame0_deriv1);
$readmemb("size12_type1_frame0_deriv2.mem", size12_type1_frame0_deriv2);
$readmemb("size12_type1_frame0_deriv3.mem", size12_type1_frame0_deriv3);
$readmemb("size12_type1_frame1_deriv0.mem", size12_type1_frame1_deriv0);
$readmemb("size12_type1_frame1_deriv1.mem", size12_type1_frame1_deriv1);
$readmemb("size12_type1_frame1_deriv2.mem", size12_type1_frame1_deriv2);
$readmemb("size12_type1_frame1_deriv3.mem", size12_type1_frame1_deriv3);
$readmemb("size13_type0_frame0_deriv0.mem", size13_type0_frame0_deriv0);
$readmemb("size13_type0_frame0_deriv1.mem", size13_type0_frame0_deriv1);
$readmemb("size13_type0_frame0_deriv2.mem", size13_type0_frame0_deriv2);
$readmemb("size13_type0_frame0_deriv3.mem", size13_type0_frame0_deriv3);
$readmemb("size13_type0_frame1_deriv0.mem", size13_type0_frame1_deriv0);
$readmemb("size13_type0_frame1_deriv1.mem", size13_type0_frame1_deriv1);
$readmemb("size13_type0_frame1_deriv2.mem", size13_type0_frame1_deriv2);
$readmemb("size13_type0_frame1_deriv3.mem", size13_type0_frame1_deriv3);
$readmemb("size13_type1_frame0_deriv0.mem", size13_type1_frame0_deriv0);
$readmemb("size13_type1_frame0_deriv1.mem", size13_type1_frame0_deriv1);
$readmemb("size13_type1_frame0_deriv2.mem", size13_type1_frame0_deriv2);
$readmemb("size13_type1_frame0_deriv3.mem", size13_type1_frame0_deriv3);
$readmemb("size13_type1_frame1_deriv0.mem", size13_type1_frame1_deriv0);
$readmemb("size13_type1_frame1_deriv1.mem", size13_type1_frame1_deriv1);
$readmemb("size13_type1_frame1_deriv2.mem", size13_type1_frame1_deriv2);
$readmemb("size13_type1_frame1_deriv3.mem", size13_type1_frame1_deriv3);
$readmemb("size14_type0_frame0_deriv0.mem", size14_type0_frame0_deriv0);
$readmemb("size14_type0_frame0_deriv1.mem", size14_type0_frame0_deriv1);
$readmemb("size14_type0_frame0_deriv2.mem", size14_type0_frame0_deriv2);
$readmemb("size14_type0_frame0_deriv3.mem", size14_type0_frame0_deriv3);
$readmemb("size14_type0_frame1_deriv0.mem", size14_type0_frame1_deriv0);
$readmemb("size14_type0_frame1_deriv1.mem", size14_type0_frame1_deriv1);
$readmemb("size14_type0_frame1_deriv2.mem", size14_type0_frame1_deriv2);
$readmemb("size14_type0_frame1_deriv3.mem", size14_type0_frame1_deriv3);
$readmemb("size14_type1_frame0_deriv0.mem", size14_type1_frame0_deriv0);
$readmemb("size14_type1_frame0_deriv1.mem", size14_type1_frame0_deriv1);
$readmemb("size14_type1_frame0_deriv2.mem", size14_type1_frame0_deriv2);
$readmemb("size14_type1_frame0_deriv3.mem", size14_type1_frame0_deriv3);
$readmemb("size14_type1_frame1_deriv0.mem", size14_type1_frame1_deriv0);
$readmemb("size14_type1_frame1_deriv1.mem", size14_type1_frame1_deriv1);
$readmemb("size14_type1_frame1_deriv2.mem", size14_type1_frame1_deriv2);
$readmemb("size14_type1_frame1_deriv3.mem", size14_type1_frame1_deriv3);
$readmemb("size15_type0_frame0_deriv0.mem", size15_type0_frame0_deriv0);
$readmemb("size15_type0_frame0_deriv1.mem", size15_type0_frame0_deriv1);
$readmemb("size15_type0_frame0_deriv2.mem", size15_type0_frame0_deriv2);
$readmemb("size15_type0_frame0_deriv3.mem", size15_type0_frame0_deriv3);
$readmemb("size15_type0_frame1_deriv0.mem", size15_type0_frame1_deriv0);
$readmemb("size15_type0_frame1_deriv1.mem", size15_type0_frame1_deriv1);
$readmemb("size15_type0_frame1_deriv2.mem", size15_type0_frame1_deriv2);
$readmemb("size15_type0_frame1_deriv3.mem", size15_type0_frame1_deriv3);
$readmemb("size15_type1_frame0_deriv0.mem", size15_type1_frame0_deriv0);
$readmemb("size15_type1_frame0_deriv1.mem", size15_type1_frame0_deriv1);
$readmemb("size15_type1_frame0_deriv2.mem", size15_type1_frame0_deriv2);
$readmemb("size15_type1_frame0_deriv3.mem", size15_type1_frame0_deriv3);
$readmemb("size15_type1_frame1_deriv0.mem", size15_type1_frame1_deriv0);
$readmemb("size15_type1_frame1_deriv1.mem", size15_type1_frame1_deriv1);
$readmemb("size15_type1_frame1_deriv2.mem", size15_type1_frame1_deriv2);
$readmemb("size15_type1_frame1_deriv3.mem", size15_type1_frame1_deriv3);
end

always @* begin
case({size_select, alien_type[1], frame_num, deriv_select})
9'b000000000: palette_out = size0_type0_frame0_deriv0[pixel_addr];
9'b000000001: palette_out = size0_type0_frame0_deriv1[pixel_addr];
9'b000000010: palette_out = size0_type0_frame0_deriv2[pixel_addr];
9'b000000011: palette_out = size0_type0_frame0_deriv3[pixel_addr];
9'b000000100: palette_out = size0_type0_frame1_deriv0[pixel_addr];
9'b000000101: palette_out = size0_type0_frame1_deriv1[pixel_addr];
9'b000000110: palette_out = size0_type0_frame1_deriv2[pixel_addr];
9'b000000111: palette_out = size0_type0_frame1_deriv3[pixel_addr];
9'b000010000: palette_out = size0_type1_frame0_deriv0[pixel_addr];
9'b000010001: palette_out = size0_type1_frame0_deriv1[pixel_addr];
9'b000010010: palette_out = size0_type1_frame0_deriv2[pixel_addr];
9'b000010011: palette_out = size0_type1_frame0_deriv3[pixel_addr];
9'b000010100: palette_out = size0_type1_frame1_deriv0[pixel_addr];
9'b000010101: palette_out = size0_type1_frame1_deriv1[pixel_addr];
9'b000010110: palette_out = size0_type1_frame1_deriv2[pixel_addr];
9'b000010111: palette_out = size0_type1_frame1_deriv3[pixel_addr];
9'b000100000: palette_out = size1_type0_frame0_deriv0[pixel_addr];
9'b000100001: palette_out = size1_type0_frame0_deriv1[pixel_addr];
9'b000100010: palette_out = size1_type0_frame0_deriv2[pixel_addr];
9'b000100011: palette_out = size1_type0_frame0_deriv3[pixel_addr];
9'b000100100: palette_out = size1_type0_frame1_deriv0[pixel_addr];
9'b000100101: palette_out = size1_type0_frame1_deriv1[pixel_addr];
9'b000100110: palette_out = size1_type0_frame1_deriv2[pixel_addr];
9'b000100111: palette_out = size1_type0_frame1_deriv3[pixel_addr];
9'b000110000: palette_out = size1_type1_frame0_deriv0[pixel_addr];
9'b000110001: palette_out = size1_type1_frame0_deriv1[pixel_addr];
9'b000110010: palette_out = size1_type1_frame0_deriv2[pixel_addr];
9'b000110011: palette_out = size1_type1_frame0_deriv3[pixel_addr];
9'b000110100: palette_out = size1_type1_frame1_deriv0[pixel_addr];
9'b000110101: palette_out = size1_type1_frame1_deriv1[pixel_addr];
9'b000110110: palette_out = size1_type1_frame1_deriv2[pixel_addr];
9'b000110111: palette_out = size1_type1_frame1_deriv3[pixel_addr];
9'b001000000: palette_out = size2_type0_frame0_deriv0[pixel_addr];
9'b001000001: palette_out = size2_type0_frame0_deriv1[pixel_addr];
9'b001000010: palette_out = size2_type0_frame0_deriv2[pixel_addr];
9'b001000011: palette_out = size2_type0_frame0_deriv3[pixel_addr];
9'b001000100: palette_out = size2_type0_frame1_deriv0[pixel_addr];
9'b001000101: palette_out = size2_type0_frame1_deriv1[pixel_addr];
9'b001000110: palette_out = size2_type0_frame1_deriv2[pixel_addr];
9'b001000111: palette_out = size2_type0_frame1_deriv3[pixel_addr];
9'b001010000: palette_out = size2_type1_frame0_deriv0[pixel_addr];
9'b001010001: palette_out = size2_type1_frame0_deriv1[pixel_addr];
9'b001010010: palette_out = size2_type1_frame0_deriv2[pixel_addr];
9'b001010011: palette_out = size2_type1_frame0_deriv3[pixel_addr];
9'b001010100: palette_out = size2_type1_frame1_deriv0[pixel_addr];
9'b001010101: palette_out = size2_type1_frame1_deriv1[pixel_addr];
9'b001010110: palette_out = size2_type1_frame1_deriv2[pixel_addr];
9'b001010111: palette_out = size2_type1_frame1_deriv3[pixel_addr];
9'b001100000: palette_out = size3_type0_frame0_deriv0[pixel_addr];
9'b001100001: palette_out = size3_type0_frame0_deriv1[pixel_addr];
9'b001100010: palette_out = size3_type0_frame0_deriv2[pixel_addr];
9'b001100011: palette_out = size3_type0_frame0_deriv3[pixel_addr];
9'b001100100: palette_out = size3_type0_frame1_deriv0[pixel_addr];
9'b001100101: palette_out = size3_type0_frame1_deriv1[pixel_addr];
9'b001100110: palette_out = size3_type0_frame1_deriv2[pixel_addr];
9'b001100111: palette_out = size3_type0_frame1_deriv3[pixel_addr];
9'b001110000: palette_out = size3_type1_frame0_deriv0[pixel_addr];
9'b001110001: palette_out = size3_type1_frame0_deriv1[pixel_addr];
9'b001110010: palette_out = size3_type1_frame0_deriv2[pixel_addr];
9'b001110011: palette_out = size3_type1_frame0_deriv3[pixel_addr];
9'b001110100: palette_out = size3_type1_frame1_deriv0[pixel_addr];
9'b001110101: palette_out = size3_type1_frame1_deriv1[pixel_addr];
9'b001110110: palette_out = size3_type1_frame1_deriv2[pixel_addr];
9'b001110111: palette_out = size3_type1_frame1_deriv3[pixel_addr];
9'b010000000: palette_out = size4_type0_frame0_deriv0[pixel_addr];
9'b010000001: palette_out = size4_type0_frame0_deriv1[pixel_addr];
9'b010000010: palette_out = size4_type0_frame0_deriv2[pixel_addr];
9'b010000011: palette_out = size4_type0_frame0_deriv3[pixel_addr];
9'b010000100: palette_out = size4_type0_frame1_deriv0[pixel_addr];
9'b010000101: palette_out = size4_type0_frame1_deriv1[pixel_addr];
9'b010000110: palette_out = size4_type0_frame1_deriv2[pixel_addr];
9'b010000111: palette_out = size4_type0_frame1_deriv3[pixel_addr];
9'b010010000: palette_out = size4_type1_frame0_deriv0[pixel_addr];
9'b010010001: palette_out = size4_type1_frame0_deriv1[pixel_addr];
9'b010010010: palette_out = size4_type1_frame0_deriv2[pixel_addr];
9'b010010011: palette_out = size4_type1_frame0_deriv3[pixel_addr];
9'b010010100: palette_out = size4_type1_frame1_deriv0[pixel_addr];
9'b010010101: palette_out = size4_type1_frame1_deriv1[pixel_addr];
9'b010010110: palette_out = size4_type1_frame1_deriv2[pixel_addr];
9'b010010111: palette_out = size4_type1_frame1_deriv3[pixel_addr];
9'b010100000: palette_out = size5_type0_frame0_deriv0[pixel_addr];
9'b010100001: palette_out = size5_type0_frame0_deriv1[pixel_addr];
9'b010100010: palette_out = size5_type0_frame0_deriv2[pixel_addr];
9'b010100011: palette_out = size5_type0_frame0_deriv3[pixel_addr];
9'b010100100: palette_out = size5_type0_frame1_deriv0[pixel_addr];
9'b010100101: palette_out = size5_type0_frame1_deriv1[pixel_addr];
9'b010100110: palette_out = size5_type0_frame1_deriv2[pixel_addr];
9'b010100111: palette_out = size5_type0_frame1_deriv3[pixel_addr];
9'b010110000: palette_out = size5_type1_frame0_deriv0[pixel_addr];
9'b010110001: palette_out = size5_type1_frame0_deriv1[pixel_addr];
9'b010110010: palette_out = size5_type1_frame0_deriv2[pixel_addr];
9'b010110011: palette_out = size5_type1_frame0_deriv3[pixel_addr];
9'b010110100: palette_out = size5_type1_frame1_deriv0[pixel_addr];
9'b010110101: palette_out = size5_type1_frame1_deriv1[pixel_addr];
9'b010110110: palette_out = size5_type1_frame1_deriv2[pixel_addr];
9'b010110111: palette_out = size5_type1_frame1_deriv3[pixel_addr];
9'b011000000: palette_out = size6_type0_frame0_deriv0[pixel_addr];
9'b011000001: palette_out = size6_type0_frame0_deriv1[pixel_addr];
9'b011000010: palette_out = size6_type0_frame0_deriv2[pixel_addr];
9'b011000011: palette_out = size6_type0_frame0_deriv3[pixel_addr];
9'b011000100: palette_out = size6_type0_frame1_deriv0[pixel_addr];
9'b011000101: palette_out = size6_type0_frame1_deriv1[pixel_addr];
9'b011000110: palette_out = size6_type0_frame1_deriv2[pixel_addr];
9'b011000111: palette_out = size6_type0_frame1_deriv3[pixel_addr];
9'b011010000: palette_out = size6_type1_frame0_deriv0[pixel_addr];
9'b011010001: palette_out = size6_type1_frame0_deriv1[pixel_addr];
9'b011010010: palette_out = size6_type1_frame0_deriv2[pixel_addr];
9'b011010011: palette_out = size6_type1_frame0_deriv3[pixel_addr];
9'b011010100: palette_out = size6_type1_frame1_deriv0[pixel_addr];
9'b011010101: palette_out = size6_type1_frame1_deriv1[pixel_addr];
9'b011010110: palette_out = size6_type1_frame1_deriv2[pixel_addr];
9'b011010111: palette_out = size6_type1_frame1_deriv3[pixel_addr];
9'b011100000: palette_out = size7_type0_frame0_deriv0[pixel_addr];
9'b011100001: palette_out = size7_type0_frame0_deriv1[pixel_addr];
9'b011100010: palette_out = size7_type0_frame0_deriv2[pixel_addr];
9'b011100011: palette_out = size7_type0_frame0_deriv3[pixel_addr];
9'b011100100: palette_out = size7_type0_frame1_deriv0[pixel_addr];
9'b011100101: palette_out = size7_type0_frame1_deriv1[pixel_addr];
9'b011100110: palette_out = size7_type0_frame1_deriv2[pixel_addr];
9'b011100111: palette_out = size7_type0_frame1_deriv3[pixel_addr];
9'b011110000: palette_out = size7_type1_frame0_deriv0[pixel_addr];
9'b011110001: palette_out = size7_type1_frame0_deriv1[pixel_addr];
9'b011110010: palette_out = size7_type1_frame0_deriv2[pixel_addr];
9'b011110011: palette_out = size7_type1_frame0_deriv3[pixel_addr];
9'b011110100: palette_out = size7_type1_frame1_deriv0[pixel_addr];
9'b011110101: palette_out = size7_type1_frame1_deriv1[pixel_addr];
9'b011110110: palette_out = size7_type1_frame1_deriv2[pixel_addr];
9'b011110111: palette_out = size7_type1_frame1_deriv3[pixel_addr];
9'b100000000: palette_out = size8_type0_frame0_deriv0[pixel_addr];
9'b100000001: palette_out = size8_type0_frame0_deriv1[pixel_addr];
9'b100000010: palette_out = size8_type0_frame0_deriv2[pixel_addr];
9'b100000011: palette_out = size8_type0_frame0_deriv3[pixel_addr];
9'b100000100: palette_out = size8_type0_frame1_deriv0[pixel_addr];
9'b100000101: palette_out = size8_type0_frame1_deriv1[pixel_addr];
9'b100000110: palette_out = size8_type0_frame1_deriv2[pixel_addr];
9'b100000111: palette_out = size8_type0_frame1_deriv3[pixel_addr];
9'b100010000: palette_out = size8_type1_frame0_deriv0[pixel_addr];
9'b100010001: palette_out = size8_type1_frame0_deriv1[pixel_addr];
9'b100010010: palette_out = size8_type1_frame0_deriv2[pixel_addr];
9'b100010011: palette_out = size8_type1_frame0_deriv3[pixel_addr];
9'b100010100: palette_out = size8_type1_frame1_deriv0[pixel_addr];
9'b100010101: palette_out = size8_type1_frame1_deriv1[pixel_addr];
9'b100010110: palette_out = size8_type1_frame1_deriv2[pixel_addr];
9'b100010111: palette_out = size8_type1_frame1_deriv3[pixel_addr];
9'b100100000: palette_out = size9_type0_frame0_deriv0[pixel_addr];
9'b100100001: palette_out = size9_type0_frame0_deriv1[pixel_addr];
9'b100100010: palette_out = size9_type0_frame0_deriv2[pixel_addr];
9'b100100011: palette_out = size9_type0_frame0_deriv3[pixel_addr];
9'b100100100: palette_out = size9_type0_frame1_deriv0[pixel_addr];
9'b100100101: palette_out = size9_type0_frame1_deriv1[pixel_addr];
9'b100100110: palette_out = size9_type0_frame1_deriv2[pixel_addr];
9'b100100111: palette_out = size9_type0_frame1_deriv3[pixel_addr];
9'b100110000: palette_out = size9_type1_frame0_deriv0[pixel_addr];
9'b100110001: palette_out = size9_type1_frame0_deriv1[pixel_addr];
9'b100110010: palette_out = size9_type1_frame0_deriv2[pixel_addr];
9'b100110011: palette_out = size9_type1_frame0_deriv3[pixel_addr];
9'b100110100: palette_out = size9_type1_frame1_deriv0[pixel_addr];
9'b100110101: palette_out = size9_type1_frame1_deriv1[pixel_addr];
9'b100110110: palette_out = size9_type1_frame1_deriv2[pixel_addr];
9'b100110111: palette_out = size9_type1_frame1_deriv3[pixel_addr];
9'b101000000: palette_out = size10_type0_frame0_deriv0[pixel_addr];
9'b101000001: palette_out = size10_type0_frame0_deriv1[pixel_addr];
9'b101000010: palette_out = size10_type0_frame0_deriv2[pixel_addr];
9'b101000011: palette_out = size10_type0_frame0_deriv3[pixel_addr];
9'b101000100: palette_out = size10_type0_frame1_deriv0[pixel_addr];
9'b101000101: palette_out = size10_type0_frame1_deriv1[pixel_addr];
9'b101000110: palette_out = size10_type0_frame1_deriv2[pixel_addr];
9'b101000111: palette_out = size10_type0_frame1_deriv3[pixel_addr];
9'b101010000: palette_out = size10_type1_frame0_deriv0[pixel_addr];
9'b101010001: palette_out = size10_type1_frame0_deriv1[pixel_addr];
9'b101010010: palette_out = size10_type1_frame0_deriv2[pixel_addr];
9'b101010011: palette_out = size10_type1_frame0_deriv3[pixel_addr];
9'b101010100: palette_out = size10_type1_frame1_deriv0[pixel_addr];
9'b101010101: palette_out = size10_type1_frame1_deriv1[pixel_addr];
9'b101010110: palette_out = size10_type1_frame1_deriv2[pixel_addr];
9'b101010111: palette_out = size10_type1_frame1_deriv3[pixel_addr];
9'b101100000: palette_out = size11_type0_frame0_deriv0[pixel_addr];
9'b101100001: palette_out = size11_type0_frame0_deriv1[pixel_addr];
9'b101100010: palette_out = size11_type0_frame0_deriv2[pixel_addr];
9'b101100011: palette_out = size11_type0_frame0_deriv3[pixel_addr];
9'b101100100: palette_out = size11_type0_frame1_deriv0[pixel_addr];
9'b101100101: palette_out = size11_type0_frame1_deriv1[pixel_addr];
9'b101100110: palette_out = size11_type0_frame1_deriv2[pixel_addr];
9'b101100111: palette_out = size11_type0_frame1_deriv3[pixel_addr];
9'b101110000: palette_out = size11_type1_frame0_deriv0[pixel_addr];
9'b101110001: palette_out = size11_type1_frame0_deriv1[pixel_addr];
9'b101110010: palette_out = size11_type1_frame0_deriv2[pixel_addr];
9'b101110011: palette_out = size11_type1_frame0_deriv3[pixel_addr];
9'b101110100: palette_out = size11_type1_frame1_deriv0[pixel_addr];
9'b101110101: palette_out = size11_type1_frame1_deriv1[pixel_addr];
9'b101110110: palette_out = size11_type1_frame1_deriv2[pixel_addr];
9'b101110111: palette_out = size11_type1_frame1_deriv3[pixel_addr];
9'b110000000: palette_out = size12_type0_frame0_deriv0[pixel_addr];
9'b110000001: palette_out = size12_type0_frame0_deriv1[pixel_addr];
9'b110000010: palette_out = size12_type0_frame0_deriv2[pixel_addr];
9'b110000011: palette_out = size12_type0_frame0_deriv3[pixel_addr];
9'b110000100: palette_out = size12_type0_frame1_deriv0[pixel_addr];
9'b110000101: palette_out = size12_type0_frame1_deriv1[pixel_addr];
9'b110000110: palette_out = size12_type0_frame1_deriv2[pixel_addr];
9'b110000111: palette_out = size12_type0_frame1_deriv3[pixel_addr];
9'b110010000: palette_out = size12_type1_frame0_deriv0[pixel_addr];
9'b110010001: palette_out = size12_type1_frame0_deriv1[pixel_addr];
9'b110010010: palette_out = size12_type1_frame0_deriv2[pixel_addr];
9'b110010011: palette_out = size12_type1_frame0_deriv3[pixel_addr];
9'b110010100: palette_out = size12_type1_frame1_deriv0[pixel_addr];
9'b110010101: palette_out = size12_type1_frame1_deriv1[pixel_addr];
9'b110010110: palette_out = size12_type1_frame1_deriv2[pixel_addr];
9'b110010111: palette_out = size12_type1_frame1_deriv3[pixel_addr];
9'b110100000: palette_out = size13_type0_frame0_deriv0[pixel_addr];
9'b110100001: palette_out = size13_type0_frame0_deriv1[pixel_addr];
9'b110100010: palette_out = size13_type0_frame0_deriv2[pixel_addr];
9'b110100011: palette_out = size13_type0_frame0_deriv3[pixel_addr];
9'b110100100: palette_out = size13_type0_frame1_deriv0[pixel_addr];
9'b110100101: palette_out = size13_type0_frame1_deriv1[pixel_addr];
9'b110100110: palette_out = size13_type0_frame1_deriv2[pixel_addr];
9'b110100111: palette_out = size13_type0_frame1_deriv3[pixel_addr];
9'b110110000: palette_out = size13_type1_frame0_deriv0[pixel_addr];
9'b110110001: palette_out = size13_type1_frame0_deriv1[pixel_addr];
9'b110110010: palette_out = size13_type1_frame0_deriv2[pixel_addr];
9'b110110011: palette_out = size13_type1_frame0_deriv3[pixel_addr];
9'b110110100: palette_out = size13_type1_frame1_deriv0[pixel_addr];
9'b110110101: palette_out = size13_type1_frame1_deriv1[pixel_addr];
9'b110110110: palette_out = size13_type1_frame1_deriv2[pixel_addr];
9'b110110111: palette_out = size13_type1_frame1_deriv3[pixel_addr];
9'b111000000: palette_out = size14_type0_frame0_deriv0[pixel_addr];
9'b111000001: palette_out = size14_type0_frame0_deriv1[pixel_addr];
9'b111000010: palette_out = size14_type0_frame0_deriv2[pixel_addr];
9'b111000011: palette_out = size14_type0_frame0_deriv3[pixel_addr];
9'b111000100: palette_out = size14_type0_frame1_deriv0[pixel_addr];
9'b111000101: palette_out = size14_type0_frame1_deriv1[pixel_addr];
9'b111000110: palette_out = size14_type0_frame1_deriv2[pixel_addr];
9'b111000111: palette_out = size14_type0_frame1_deriv3[pixel_addr];
9'b111010000: palette_out = size14_type1_frame0_deriv0[pixel_addr];
9'b111010001: palette_out = size14_type1_frame0_deriv1[pixel_addr];
9'b111010010: palette_out = size14_type1_frame0_deriv2[pixel_addr];
9'b111010011: palette_out = size14_type1_frame0_deriv3[pixel_addr];
9'b111010100: palette_out = size14_type1_frame1_deriv0[pixel_addr];
9'b111010101: palette_out = size14_type1_frame1_deriv1[pixel_addr];
9'b111010110: palette_out = size14_type1_frame1_deriv2[pixel_addr];
9'b111010111: palette_out = size14_type1_frame1_deriv3[pixel_addr];
9'b111100000: palette_out = size15_type0_frame0_deriv0[pixel_addr];
9'b111100001: palette_out = size15_type0_frame0_deriv1[pixel_addr];
9'b111100010: palette_out = size15_type0_frame0_deriv2[pixel_addr];
9'b111100011: palette_out = size15_type0_frame0_deriv3[pixel_addr];
9'b111100100: palette_out = size15_type0_frame1_deriv0[pixel_addr];
9'b111100101: palette_out = size15_type0_frame1_deriv1[pixel_addr];
9'b111100110: palette_out = size15_type0_frame1_deriv2[pixel_addr];
9'b111100111: palette_out = size15_type0_frame1_deriv3[pixel_addr];
9'b111110000: palette_out = size15_type1_frame0_deriv0[pixel_addr];
9'b111110001: palette_out = size15_type1_frame0_deriv1[pixel_addr];
9'b111110010: palette_out = size15_type1_frame0_deriv2[pixel_addr];
9'b111110011: palette_out = size15_type1_frame0_deriv3[pixel_addr];
9'b111110100: palette_out = size15_type1_frame1_deriv0[pixel_addr];
9'b111110101: palette_out = size15_type1_frame1_deriv1[pixel_addr];
9'b111110110: palette_out = size15_type1_frame1_deriv2[pixel_addr];
9'b111110111: palette_out = size15_type1_frame1_deriv3[pixel_addr];
default : palette_out = 0;
endcase
end
endmodule

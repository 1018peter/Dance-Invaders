`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/01/02 13:57:31
// Design Name: 
// Module Name: alien_pixel_reader
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module alien_pixel_reader(
    input [1:0] frame_num,
    input [1:0] alien_type,
    input [3:0] size_select,
    input [1:0] deriv_select,
    input [15:0] pixel_addr,
    output logic palette_out
    );
    
    
reg size0_type0_frame0_deriv0 [0:2047];
reg size0_type0_frame0_deriv1 [0:2047];
reg size0_type0_frame0_deriv2 [0:2047];
reg size0_type0_frame0_deriv3 [0:2047];
reg size0_type0_frame1_deriv0 [0:2047];
reg size0_type0_frame1_deriv1 [0:2047];
reg size0_type0_frame1_deriv2 [0:2047];
reg size0_type0_frame1_deriv3 [0:2047];
reg size0_type1_frame0_deriv0 [0:2047];
reg size0_type1_frame0_deriv1 [0:2047];
reg size0_type1_frame0_deriv2 [0:2047];
reg size0_type1_frame0_deriv3 [0:2047];
reg size0_type1_frame1_deriv0 [0:2047];
reg size0_type1_frame1_deriv1 [0:2047];
reg size0_type1_frame1_deriv2 [0:2047];
reg size0_type1_frame1_deriv3 [0:2047];
reg size1_type0_frame0_deriv0 [0:1921];
reg size1_type0_frame0_deriv1 [0:1921];
reg size1_type0_frame0_deriv2 [0:1921];
reg size1_type0_frame0_deriv3 [0:1921];
reg size1_type0_frame1_deriv0 [0:1921];
reg size1_type0_frame1_deriv1 [0:1921];
reg size1_type0_frame1_deriv2 [0:1921];
reg size1_type0_frame1_deriv3 [0:1921];
reg size1_type1_frame0_deriv0 [0:1921];
reg size1_type1_frame0_deriv1 [0:1921];
reg size1_type1_frame0_deriv2 [0:1921];
reg size1_type1_frame0_deriv3 [0:1921];
reg size1_type1_frame1_deriv0 [0:1921];
reg size1_type1_frame1_deriv1 [0:1921];
reg size1_type1_frame1_deriv2 [0:1921];
reg size1_type1_frame1_deriv3 [0:1921];
reg size2_type0_frame0_deriv0 [0:1799];
reg size2_type0_frame0_deriv1 [0:1799];
reg size2_type0_frame0_deriv2 [0:1799];
reg size2_type0_frame0_deriv3 [0:1799];
reg size2_type0_frame1_deriv0 [0:1799];
reg size2_type0_frame1_deriv1 [0:1799];
reg size2_type0_frame1_deriv2 [0:1799];
reg size2_type0_frame1_deriv3 [0:1799];
reg size2_type1_frame0_deriv0 [0:1799];
reg size2_type1_frame0_deriv1 [0:1799];
reg size2_type1_frame0_deriv2 [0:1799];
reg size2_type1_frame0_deriv3 [0:1799];
reg size2_type1_frame1_deriv0 [0:1799];
reg size2_type1_frame1_deriv1 [0:1799];
reg size2_type1_frame1_deriv2 [0:1799];
reg size2_type1_frame1_deriv3 [0:1799];
reg size3_type0_frame0_deriv0 [0:1681];
reg size3_type0_frame0_deriv1 [0:1681];
reg size3_type0_frame0_deriv2 [0:1681];
reg size3_type0_frame0_deriv3 [0:1681];
reg size3_type0_frame1_deriv0 [0:1681];
reg size3_type0_frame1_deriv1 [0:1681];
reg size3_type0_frame1_deriv2 [0:1681];
reg size3_type0_frame1_deriv3 [0:1681];
reg size3_type1_frame0_deriv0 [0:1681];
reg size3_type1_frame0_deriv1 [0:1681];
reg size3_type1_frame0_deriv2 [0:1681];
reg size3_type1_frame0_deriv3 [0:1681];
reg size3_type1_frame1_deriv0 [0:1681];
reg size3_type1_frame1_deriv1 [0:1681];
reg size3_type1_frame1_deriv2 [0:1681];
reg size3_type1_frame1_deriv3 [0:1681];
reg size4_type0_frame0_deriv0 [0:1567];
reg size4_type0_frame0_deriv1 [0:1567];
reg size4_type0_frame0_deriv2 [0:1567];
reg size4_type0_frame0_deriv3 [0:1567];
reg size4_type0_frame1_deriv0 [0:1567];
reg size4_type0_frame1_deriv1 [0:1567];
reg size4_type0_frame1_deriv2 [0:1567];
reg size4_type0_frame1_deriv3 [0:1567];
reg size4_type1_frame0_deriv0 [0:1567];
reg size4_type1_frame0_deriv1 [0:1567];
reg size4_type1_frame0_deriv2 [0:1567];
reg size4_type1_frame0_deriv3 [0:1567];
reg size4_type1_frame1_deriv0 [0:1567];
reg size4_type1_frame1_deriv1 [0:1567];
reg size4_type1_frame1_deriv2 [0:1567];
reg size4_type1_frame1_deriv3 [0:1567];
reg size5_type0_frame0_deriv0 [0:1457];
reg size5_type0_frame0_deriv1 [0:1457];
reg size5_type0_frame0_deriv2 [0:1457];
reg size5_type0_frame0_deriv3 [0:1457];
reg size5_type0_frame1_deriv0 [0:1457];
reg size5_type0_frame1_deriv1 [0:1457];
reg size5_type0_frame1_deriv2 [0:1457];
reg size5_type0_frame1_deriv3 [0:1457];
reg size5_type1_frame0_deriv0 [0:1457];
reg size5_type1_frame0_deriv1 [0:1457];
reg size5_type1_frame0_deriv2 [0:1457];
reg size5_type1_frame0_deriv3 [0:1457];
reg size5_type1_frame1_deriv0 [0:1457];
reg size5_type1_frame1_deriv1 [0:1457];
reg size5_type1_frame1_deriv2 [0:1457];
reg size5_type1_frame1_deriv3 [0:1457];
reg size6_type0_frame0_deriv0 [0:1351];
reg size6_type0_frame0_deriv1 [0:1351];
reg size6_type0_frame0_deriv2 [0:1351];
reg size6_type0_frame0_deriv3 [0:1351];
reg size6_type0_frame1_deriv0 [0:1351];
reg size6_type0_frame1_deriv1 [0:1351];
reg size6_type0_frame1_deriv2 [0:1351];
reg size6_type0_frame1_deriv3 [0:1351];
reg size6_type1_frame0_deriv0 [0:1351];
reg size6_type1_frame0_deriv1 [0:1351];
reg size6_type1_frame0_deriv2 [0:1351];
reg size6_type1_frame0_deriv3 [0:1351];
reg size6_type1_frame1_deriv0 [0:1351];
reg size6_type1_frame1_deriv1 [0:1351];
reg size6_type1_frame1_deriv2 [0:1351];
reg size6_type1_frame1_deriv3 [0:1351];
reg size7_type0_frame0_deriv0 [0:1249];
reg size7_type0_frame0_deriv1 [0:1249];
reg size7_type0_frame0_deriv2 [0:1249];
reg size7_type0_frame0_deriv3 [0:1249];
reg size7_type0_frame1_deriv0 [0:1249];
reg size7_type0_frame1_deriv1 [0:1249];
reg size7_type0_frame1_deriv2 [0:1249];
reg size7_type0_frame1_deriv3 [0:1249];
reg size7_type1_frame0_deriv0 [0:1249];
reg size7_type1_frame0_deriv1 [0:1249];
reg size7_type1_frame0_deriv2 [0:1249];
reg size7_type1_frame0_deriv3 [0:1249];
reg size7_type1_frame1_deriv0 [0:1249];
reg size7_type1_frame1_deriv1 [0:1249];
reg size7_type1_frame1_deriv2 [0:1249];
reg size7_type1_frame1_deriv3 [0:1249];
reg size8_type0_frame0_deriv0 [0:1151];
reg size8_type0_frame0_deriv1 [0:1151];
reg size8_type0_frame0_deriv2 [0:1151];
reg size8_type0_frame0_deriv3 [0:1151];
reg size8_type0_frame1_deriv0 [0:1151];
reg size8_type0_frame1_deriv1 [0:1151];
reg size8_type0_frame1_deriv2 [0:1151];
reg size8_type0_frame1_deriv3 [0:1151];
reg size8_type1_frame0_deriv0 [0:1151];
reg size8_type1_frame0_deriv1 [0:1151];
reg size8_type1_frame0_deriv2 [0:1151];
reg size8_type1_frame0_deriv3 [0:1151];
reg size8_type1_frame1_deriv0 [0:1151];
reg size8_type1_frame1_deriv1 [0:1151];
reg size8_type1_frame1_deriv2 [0:1151];
reg size8_type1_frame1_deriv3 [0:1151];
reg size9_type0_frame0_deriv0 [0:1057];
reg size9_type0_frame0_deriv1 [0:1057];
reg size9_type0_frame0_deriv2 [0:1057];
reg size9_type0_frame0_deriv3 [0:1057];
reg size9_type0_frame1_deriv0 [0:1057];
reg size9_type0_frame1_deriv1 [0:1057];
reg size9_type0_frame1_deriv2 [0:1057];
reg size9_type0_frame1_deriv3 [0:1057];
reg size9_type1_frame0_deriv0 [0:1057];
reg size9_type1_frame0_deriv1 [0:1057];
reg size9_type1_frame0_deriv2 [0:1057];
reg size9_type1_frame0_deriv3 [0:1057];
reg size9_type1_frame1_deriv0 [0:1057];
reg size9_type1_frame1_deriv1 [0:1057];
reg size9_type1_frame1_deriv2 [0:1057];
reg size9_type1_frame1_deriv3 [0:1057];
reg size10_type0_frame0_deriv0 [0:967];
reg size10_type0_frame0_deriv1 [0:967];
reg size10_type0_frame0_deriv2 [0:967];
reg size10_type0_frame0_deriv3 [0:967];
reg size10_type0_frame1_deriv0 [0:967];
reg size10_type0_frame1_deriv1 [0:967];
reg size10_type0_frame1_deriv2 [0:967];
reg size10_type0_frame1_deriv3 [0:967];
reg size10_type1_frame0_deriv0 [0:967];
reg size10_type1_frame0_deriv1 [0:967];
reg size10_type1_frame0_deriv2 [0:967];
reg size10_type1_frame0_deriv3 [0:967];
reg size10_type1_frame1_deriv0 [0:967];
reg size10_type1_frame1_deriv1 [0:967];
reg size10_type1_frame1_deriv2 [0:967];
reg size10_type1_frame1_deriv3 [0:967];
reg size11_type0_frame0_deriv0 [0:881];
reg size11_type0_frame0_deriv1 [0:881];
reg size11_type0_frame0_deriv2 [0:881];
reg size11_type0_frame0_deriv3 [0:881];
reg size11_type0_frame1_deriv0 [0:881];
reg size11_type0_frame1_deriv1 [0:881];
reg size11_type0_frame1_deriv2 [0:881];
reg size11_type0_frame1_deriv3 [0:881];
reg size11_type1_frame0_deriv0 [0:881];
reg size11_type1_frame0_deriv1 [0:881];
reg size11_type1_frame0_deriv2 [0:881];
reg size11_type1_frame0_deriv3 [0:881];
reg size11_type1_frame1_deriv0 [0:881];
reg size11_type1_frame1_deriv1 [0:881];
reg size11_type1_frame1_deriv2 [0:881];
reg size11_type1_frame1_deriv3 [0:881];
reg size12_type0_frame0_deriv0 [0:799];
reg size12_type0_frame0_deriv1 [0:799];
reg size12_type0_frame0_deriv2 [0:799];
reg size12_type0_frame0_deriv3 [0:799];
reg size12_type0_frame1_deriv0 [0:799];
reg size12_type0_frame1_deriv1 [0:799];
reg size12_type0_frame1_deriv2 [0:799];
reg size12_type0_frame1_deriv3 [0:799];
reg size12_type1_frame0_deriv0 [0:799];
reg size12_type1_frame0_deriv1 [0:799];
reg size12_type1_frame0_deriv2 [0:799];
reg size12_type1_frame0_deriv3 [0:799];
reg size12_type1_frame1_deriv0 [0:799];
reg size12_type1_frame1_deriv1 [0:799];
reg size12_type1_frame1_deriv2 [0:799];
reg size12_type1_frame1_deriv3 [0:799];
reg size13_type0_frame0_deriv0 [0:721];
reg size13_type0_frame0_deriv1 [0:721];
reg size13_type0_frame0_deriv2 [0:721];
reg size13_type0_frame0_deriv3 [0:721];
reg size13_type0_frame1_deriv0 [0:721];
reg size13_type0_frame1_deriv1 [0:721];
reg size13_type0_frame1_deriv2 [0:721];
reg size13_type0_frame1_deriv3 [0:721];
reg size13_type1_frame0_deriv0 [0:721];
reg size13_type1_frame0_deriv1 [0:721];
reg size13_type1_frame0_deriv2 [0:721];
reg size13_type1_frame0_deriv3 [0:721];
reg size13_type1_frame1_deriv0 [0:721];
reg size13_type1_frame1_deriv1 [0:721];
reg size13_type1_frame1_deriv2 [0:721];
reg size13_type1_frame1_deriv3 [0:721];
reg size14_type0_frame0_deriv0 [0:647];
reg size14_type0_frame0_deriv1 [0:647];
reg size14_type0_frame0_deriv2 [0:647];
reg size14_type0_frame0_deriv3 [0:647];
reg size14_type0_frame1_deriv0 [0:647];
reg size14_type0_frame1_deriv1 [0:647];
reg size14_type0_frame1_deriv2 [0:647];
reg size14_type0_frame1_deriv3 [0:647];
reg size14_type1_frame0_deriv0 [0:647];
reg size14_type1_frame0_deriv1 [0:647];
reg size14_type1_frame0_deriv2 [0:647];
reg size14_type1_frame0_deriv3 [0:647];
reg size14_type1_frame1_deriv0 [0:647];
reg size14_type1_frame1_deriv1 [0:647];
reg size14_type1_frame1_deriv2 [0:647];
reg size14_type1_frame1_deriv3 [0:647];
reg size15_type0_frame0_deriv0 [0:577];
reg size15_type0_frame0_deriv1 [0:577];
reg size15_type0_frame0_deriv2 [0:577];
reg size15_type0_frame0_deriv3 [0:577];
reg size15_type0_frame1_deriv0 [0:577];
reg size15_type0_frame1_deriv1 [0:577];
reg size15_type0_frame1_deriv2 [0:577];
reg size15_type0_frame1_deriv3 [0:577];
reg size15_type1_frame0_deriv0 [0:577];
reg size15_type1_frame0_deriv1 [0:577];
reg size15_type1_frame0_deriv2 [0:577];
reg size15_type1_frame0_deriv3 [0:577];
reg size15_type1_frame1_deriv0 [0:577];
reg size15_type1_frame1_deriv1 [0:577];
reg size15_type1_frame1_deriv2 [0:577];
reg size15_type1_frame1_deriv3 [0:577];


initial begin
$readmemb("size0_type0_frame0_deriv0.mem", size0_type0_frame0_deriv0);
$readmemb("size0_type0_frame0_deriv1.mem", size0_type0_frame0_deriv1);
$readmemb("size0_type0_frame0_deriv2.mem", size0_type0_frame0_deriv2);
$readmemb("size0_type0_frame0_deriv3.mem", size0_type0_frame0_deriv3);
$readmemb("size0_type0_frame1_deriv0.mem", size0_type0_frame1_deriv0);
$readmemb("size0_type0_frame1_deriv1.mem", size0_type0_frame1_deriv1);
$readmemb("size0_type0_frame1_deriv2.mem", size0_type0_frame1_deriv2);
$readmemb("size0_type0_frame1_deriv3.mem", size0_type0_frame1_deriv3);
$readmemb("size0_type1_frame0_deriv0.mem", size0_type1_frame0_deriv0);
$readmemb("size0_type1_frame0_deriv1.mem", size0_type1_frame0_deriv1);
$readmemb("size0_type1_frame0_deriv2.mem", size0_type1_frame0_deriv2);
$readmemb("size0_type1_frame0_deriv3.mem", size0_type1_frame0_deriv3);
$readmemb("size0_type1_frame1_deriv0.mem", size0_type1_frame1_deriv0);
$readmemb("size0_type1_frame1_deriv1.mem", size0_type1_frame1_deriv1);
$readmemb("size0_type1_frame1_deriv2.mem", size0_type1_frame1_deriv2);
$readmemb("size0_type1_frame1_deriv3.mem", size0_type1_frame1_deriv3);
$readmemb("size1_type0_frame0_deriv0.mem", size1_type0_frame0_deriv0);
$readmemb("size1_type0_frame0_deriv1.mem", size1_type0_frame0_deriv1);
$readmemb("size1_type0_frame0_deriv2.mem", size1_type0_frame0_deriv2);
$readmemb("size1_type0_frame0_deriv3.mem", size1_type0_frame0_deriv3);
$readmemb("size1_type0_frame1_deriv0.mem", size1_type0_frame1_deriv0);
$readmemb("size1_type0_frame1_deriv1.mem", size1_type0_frame1_deriv1);
$readmemb("size1_type0_frame1_deriv2.mem", size1_type0_frame1_deriv2);
$readmemb("size1_type0_frame1_deriv3.mem", size1_type0_frame1_deriv3);
$readmemb("size1_type1_frame0_deriv0.mem", size1_type1_frame0_deriv0);
$readmemb("size1_type1_frame0_deriv1.mem", size1_type1_frame0_deriv1);
$readmemb("size1_type1_frame0_deriv2.mem", size1_type1_frame0_deriv2);
$readmemb("size1_type1_frame0_deriv3.mem", size1_type1_frame0_deriv3);
$readmemb("size1_type1_frame1_deriv0.mem", size1_type1_frame1_deriv0);
$readmemb("size1_type1_frame1_deriv1.mem", size1_type1_frame1_deriv1);
$readmemb("size1_type1_frame1_deriv2.mem", size1_type1_frame1_deriv2);
$readmemb("size1_type1_frame1_deriv3.mem", size1_type1_frame1_deriv3);
$readmemb("size2_type0_frame0_deriv0.mem", size2_type0_frame0_deriv0);
$readmemb("size2_type0_frame0_deriv1.mem", size2_type0_frame0_deriv1);
$readmemb("size2_type0_frame0_deriv2.mem", size2_type0_frame0_deriv2);
$readmemb("size2_type0_frame0_deriv3.mem", size2_type0_frame0_deriv3);
$readmemb("size2_type0_frame1_deriv0.mem", size2_type0_frame1_deriv0);
$readmemb("size2_type0_frame1_deriv1.mem", size2_type0_frame1_deriv1);
$readmemb("size2_type0_frame1_deriv2.mem", size2_type0_frame1_deriv2);
$readmemb("size2_type0_frame1_deriv3.mem", size2_type0_frame1_deriv3);
$readmemb("size2_type1_frame0_deriv0.mem", size2_type1_frame0_deriv0);
$readmemb("size2_type1_frame0_deriv1.mem", size2_type1_frame0_deriv1);
$readmemb("size2_type1_frame0_deriv2.mem", size2_type1_frame0_deriv2);
$readmemb("size2_type1_frame0_deriv3.mem", size2_type1_frame0_deriv3);
$readmemb("size2_type1_frame1_deriv0.mem", size2_type1_frame1_deriv0);
$readmemb("size2_type1_frame1_deriv1.mem", size2_type1_frame1_deriv1);
$readmemb("size2_type1_frame1_deriv2.mem", size2_type1_frame1_deriv2);
$readmemb("size2_type1_frame1_deriv3.mem", size2_type1_frame1_deriv3);
$readmemb("size3_type0_frame0_deriv0.mem", size3_type0_frame0_deriv0);
$readmemb("size3_type0_frame0_deriv1.mem", size3_type0_frame0_deriv1);
$readmemb("size3_type0_frame0_deriv2.mem", size3_type0_frame0_deriv2);
$readmemb("size3_type0_frame0_deriv3.mem", size3_type0_frame0_deriv3);
$readmemb("size3_type0_frame1_deriv0.mem", size3_type0_frame1_deriv0);
$readmemb("size3_type0_frame1_deriv1.mem", size3_type0_frame1_deriv1);
$readmemb("size3_type0_frame1_deriv2.mem", size3_type0_frame1_deriv2);
$readmemb("size3_type0_frame1_deriv3.mem", size3_type0_frame1_deriv3);
$readmemb("size3_type1_frame0_deriv0.mem", size3_type1_frame0_deriv0);
$readmemb("size3_type1_frame0_deriv1.mem", size3_type1_frame0_deriv1);
$readmemb("size3_type1_frame0_deriv2.mem", size3_type1_frame0_deriv2);
$readmemb("size3_type1_frame0_deriv3.mem", size3_type1_frame0_deriv3);
$readmemb("size3_type1_frame1_deriv0.mem", size3_type1_frame1_deriv0);
$readmemb("size3_type1_frame1_deriv1.mem", size3_type1_frame1_deriv1);
$readmemb("size3_type1_frame1_deriv2.mem", size3_type1_frame1_deriv2);
$readmemb("size3_type1_frame1_deriv3.mem", size3_type1_frame1_deriv3);
$readmemb("size4_type0_frame0_deriv0.mem", size4_type0_frame0_deriv0);
$readmemb("size4_type0_frame0_deriv1.mem", size4_type0_frame0_deriv1);
$readmemb("size4_type0_frame0_deriv2.mem", size4_type0_frame0_deriv2);
$readmemb("size4_type0_frame0_deriv3.mem", size4_type0_frame0_deriv3);
$readmemb("size4_type0_frame1_deriv0.mem", size4_type0_frame1_deriv0);
$readmemb("size4_type0_frame1_deriv1.mem", size4_type0_frame1_deriv1);
$readmemb("size4_type0_frame1_deriv2.mem", size4_type0_frame1_deriv2);
$readmemb("size4_type0_frame1_deriv3.mem", size4_type0_frame1_deriv3);
$readmemb("size4_type1_frame0_deriv0.mem", size4_type1_frame0_deriv0);
$readmemb("size4_type1_frame0_deriv1.mem", size4_type1_frame0_deriv1);
$readmemb("size4_type1_frame0_deriv2.mem", size4_type1_frame0_deriv2);
$readmemb("size4_type1_frame0_deriv3.mem", size4_type1_frame0_deriv3);
$readmemb("size4_type1_frame1_deriv0.mem", size4_type1_frame1_deriv0);
$readmemb("size4_type1_frame1_deriv1.mem", size4_type1_frame1_deriv1);
$readmemb("size4_type1_frame1_deriv2.mem", size4_type1_frame1_deriv2);
$readmemb("size4_type1_frame1_deriv3.mem", size4_type1_frame1_deriv3);
$readmemb("size5_type0_frame0_deriv0.mem", size5_type0_frame0_deriv0);
$readmemb("size5_type0_frame0_deriv1.mem", size5_type0_frame0_deriv1);
$readmemb("size5_type0_frame0_deriv2.mem", size5_type0_frame0_deriv2);
$readmemb("size5_type0_frame0_deriv3.mem", size5_type0_frame0_deriv3);
$readmemb("size5_type0_frame1_deriv0.mem", size5_type0_frame1_deriv0);
$readmemb("size5_type0_frame1_deriv1.mem", size5_type0_frame1_deriv1);
$readmemb("size5_type0_frame1_deriv2.mem", size5_type0_frame1_deriv2);
$readmemb("size5_type0_frame1_deriv3.mem", size5_type0_frame1_deriv3);
$readmemb("size5_type1_frame0_deriv0.mem", size5_type1_frame0_deriv0);
$readmemb("size5_type1_frame0_deriv1.mem", size5_type1_frame0_deriv1);
$readmemb("size5_type1_frame0_deriv2.mem", size5_type1_frame0_deriv2);
$readmemb("size5_type1_frame0_deriv3.mem", size5_type1_frame0_deriv3);
$readmemb("size5_type1_frame1_deriv0.mem", size5_type1_frame1_deriv0);
$readmemb("size5_type1_frame1_deriv1.mem", size5_type1_frame1_deriv1);
$readmemb("size5_type1_frame1_deriv2.mem", size5_type1_frame1_deriv2);
$readmemb("size5_type1_frame1_deriv3.mem", size5_type1_frame1_deriv3);
$readmemb("size6_type0_frame0_deriv0.mem", size6_type0_frame0_deriv0);
$readmemb("size6_type0_frame0_deriv1.mem", size6_type0_frame0_deriv1);
$readmemb("size6_type0_frame0_deriv2.mem", size6_type0_frame0_deriv2);
$readmemb("size6_type0_frame0_deriv3.mem", size6_type0_frame0_deriv3);
$readmemb("size6_type0_frame1_deriv0.mem", size6_type0_frame1_deriv0);
$readmemb("size6_type0_frame1_deriv1.mem", size6_type0_frame1_deriv1);
$readmemb("size6_type0_frame1_deriv2.mem", size6_type0_frame1_deriv2);
$readmemb("size6_type0_frame1_deriv3.mem", size6_type0_frame1_deriv3);
$readmemb("size6_type1_frame0_deriv0.mem", size6_type1_frame0_deriv0);
$readmemb("size6_type1_frame0_deriv1.mem", size6_type1_frame0_deriv1);
$readmemb("size6_type1_frame0_deriv2.mem", size6_type1_frame0_deriv2);
$readmemb("size6_type1_frame0_deriv3.mem", size6_type1_frame0_deriv3);
$readmemb("size6_type1_frame1_deriv0.mem", size6_type1_frame1_deriv0);
$readmemb("size6_type1_frame1_deriv1.mem", size6_type1_frame1_deriv1);
$readmemb("size6_type1_frame1_deriv2.mem", size6_type1_frame1_deriv2);
$readmemb("size6_type1_frame1_deriv3.mem", size6_type1_frame1_deriv3);
$readmemb("size7_type0_frame0_deriv0.mem", size7_type0_frame0_deriv0);
$readmemb("size7_type0_frame0_deriv1.mem", size7_type0_frame0_deriv1);
$readmemb("size7_type0_frame0_deriv2.mem", size7_type0_frame0_deriv2);
$readmemb("size7_type0_frame0_deriv3.mem", size7_type0_frame0_deriv3);
$readmemb("size7_type0_frame1_deriv0.mem", size7_type0_frame1_deriv0);
$readmemb("size7_type0_frame1_deriv1.mem", size7_type0_frame1_deriv1);
$readmemb("size7_type0_frame1_deriv2.mem", size7_type0_frame1_deriv2);
$readmemb("size7_type0_frame1_deriv3.mem", size7_type0_frame1_deriv3);
$readmemb("size7_type1_frame0_deriv0.mem", size7_type1_frame0_deriv0);
$readmemb("size7_type1_frame0_deriv1.mem", size7_type1_frame0_deriv1);
$readmemb("size7_type1_frame0_deriv2.mem", size7_type1_frame0_deriv2);
$readmemb("size7_type1_frame0_deriv3.mem", size7_type1_frame0_deriv3);
$readmemb("size7_type1_frame1_deriv0.mem", size7_type1_frame1_deriv0);
$readmemb("size7_type1_frame1_deriv1.mem", size7_type1_frame1_deriv1);
$readmemb("size7_type1_frame1_deriv2.mem", size7_type1_frame1_deriv2);
$readmemb("size7_type1_frame1_deriv3.mem", size7_type1_frame1_deriv3);
$readmemb("size8_type0_frame0_deriv0.mem", size8_type0_frame0_deriv0);
$readmemb("size8_type0_frame0_deriv1.mem", size8_type0_frame0_deriv1);
$readmemb("size8_type0_frame0_deriv2.mem", size8_type0_frame0_deriv2);
$readmemb("size8_type0_frame0_deriv3.mem", size8_type0_frame0_deriv3);
$readmemb("size8_type0_frame1_deriv0.mem", size8_type0_frame1_deriv0);
$readmemb("size8_type0_frame1_deriv1.mem", size8_type0_frame1_deriv1);
$readmemb("size8_type0_frame1_deriv2.mem", size8_type0_frame1_deriv2);
$readmemb("size8_type0_frame1_deriv3.mem", size8_type0_frame1_deriv3);
$readmemb("size8_type1_frame0_deriv0.mem", size8_type1_frame0_deriv0);
$readmemb("size8_type1_frame0_deriv1.mem", size8_type1_frame0_deriv1);
$readmemb("size8_type1_frame0_deriv2.mem", size8_type1_frame0_deriv2);
$readmemb("size8_type1_frame0_deriv3.mem", size8_type1_frame0_deriv3);
$readmemb("size8_type1_frame1_deriv0.mem", size8_type1_frame1_deriv0);
$readmemb("size8_type1_frame1_deriv1.mem", size8_type1_frame1_deriv1);
$readmemb("size8_type1_frame1_deriv2.mem", size8_type1_frame1_deriv2);
$readmemb("size8_type1_frame1_deriv3.mem", size8_type1_frame1_deriv3);
$readmemb("size9_type0_frame0_deriv0.mem", size9_type0_frame0_deriv0);
$readmemb("size9_type0_frame0_deriv1.mem", size9_type0_frame0_deriv1);
$readmemb("size9_type0_frame0_deriv2.mem", size9_type0_frame0_deriv2);
$readmemb("size9_type0_frame0_deriv3.mem", size9_type0_frame0_deriv3);
$readmemb("size9_type0_frame1_deriv0.mem", size9_type0_frame1_deriv0);
$readmemb("size9_type0_frame1_deriv1.mem", size9_type0_frame1_deriv1);
$readmemb("size9_type0_frame1_deriv2.mem", size9_type0_frame1_deriv2);
$readmemb("size9_type0_frame1_deriv3.mem", size9_type0_frame1_deriv3);
$readmemb("size9_type1_frame0_deriv0.mem", size9_type1_frame0_deriv0);
$readmemb("size9_type1_frame0_deriv1.mem", size9_type1_frame0_deriv1);
$readmemb("size9_type1_frame0_deriv2.mem", size9_type1_frame0_deriv2);
$readmemb("size9_type1_frame0_deriv3.mem", size9_type1_frame0_deriv3);
$readmemb("size9_type1_frame1_deriv0.mem", size9_type1_frame1_deriv0);
$readmemb("size9_type1_frame1_deriv1.mem", size9_type1_frame1_deriv1);
$readmemb("size9_type1_frame1_deriv2.mem", size9_type1_frame1_deriv2);
$readmemb("size9_type1_frame1_deriv3.mem", size9_type1_frame1_deriv3);
$readmemb("size10_type0_frame0_deriv0.mem", size10_type0_frame0_deriv0);
$readmemb("size10_type0_frame0_deriv1.mem", size10_type0_frame0_deriv1);
$readmemb("size10_type0_frame0_deriv2.mem", size10_type0_frame0_deriv2);
$readmemb("size10_type0_frame0_deriv3.mem", size10_type0_frame0_deriv3);
$readmemb("size10_type0_frame1_deriv0.mem", size10_type0_frame1_deriv0);
$readmemb("size10_type0_frame1_deriv1.mem", size10_type0_frame1_deriv1);
$readmemb("size10_type0_frame1_deriv2.mem", size10_type0_frame1_deriv2);
$readmemb("size10_type0_frame1_deriv3.mem", size10_type0_frame1_deriv3);
$readmemb("size10_type1_frame0_deriv0.mem", size10_type1_frame0_deriv0);
$readmemb("size10_type1_frame0_deriv1.mem", size10_type1_frame0_deriv1);
$readmemb("size10_type1_frame0_deriv2.mem", size10_type1_frame0_deriv2);
$readmemb("size10_type1_frame0_deriv3.mem", size10_type1_frame0_deriv3);
$readmemb("size10_type1_frame1_deriv0.mem", size10_type1_frame1_deriv0);
$readmemb("size10_type1_frame1_deriv1.mem", size10_type1_frame1_deriv1);
$readmemb("size10_type1_frame1_deriv2.mem", size10_type1_frame1_deriv2);
$readmemb("size10_type1_frame1_deriv3.mem", size10_type1_frame1_deriv3);
$readmemb("size11_type0_frame0_deriv0.mem", size11_type0_frame0_deriv0);
$readmemb("size11_type0_frame0_deriv1.mem", size11_type0_frame0_deriv1);
$readmemb("size11_type0_frame0_deriv2.mem", size11_type0_frame0_deriv2);
$readmemb("size11_type0_frame0_deriv3.mem", size11_type0_frame0_deriv3);
$readmemb("size11_type0_frame1_deriv0.mem", size11_type0_frame1_deriv0);
$readmemb("size11_type0_frame1_deriv1.mem", size11_type0_frame1_deriv1);
$readmemb("size11_type0_frame1_deriv2.mem", size11_type0_frame1_deriv2);
$readmemb("size11_type0_frame1_deriv3.mem", size11_type0_frame1_deriv3);
$readmemb("size11_type1_frame0_deriv0.mem", size11_type1_frame0_deriv0);
$readmemb("size11_type1_frame0_deriv1.mem", size11_type1_frame0_deriv1);
$readmemb("size11_type1_frame0_deriv2.mem", size11_type1_frame0_deriv2);
$readmemb("size11_type1_frame0_deriv3.mem", size11_type1_frame0_deriv3);
$readmemb("size11_type1_frame1_deriv0.mem", size11_type1_frame1_deriv0);
$readmemb("size11_type1_frame1_deriv1.mem", size11_type1_frame1_deriv1);
$readmemb("size11_type1_frame1_deriv2.mem", size11_type1_frame1_deriv2);
$readmemb("size11_type1_frame1_deriv3.mem", size11_type1_frame1_deriv3);
$readmemb("size12_type0_frame0_deriv0.mem", size12_type0_frame0_deriv0);
$readmemb("size12_type0_frame0_deriv1.mem", size12_type0_frame0_deriv1);
$readmemb("size12_type0_frame0_deriv2.mem", size12_type0_frame0_deriv2);
$readmemb("size12_type0_frame0_deriv3.mem", size12_type0_frame0_deriv3);
$readmemb("size12_type0_frame1_deriv0.mem", size12_type0_frame1_deriv0);
$readmemb("size12_type0_frame1_deriv1.mem", size12_type0_frame1_deriv1);
$readmemb("size12_type0_frame1_deriv2.mem", size12_type0_frame1_deriv2);
$readmemb("size12_type0_frame1_deriv3.mem", size12_type0_frame1_deriv3);
$readmemb("size12_type1_frame0_deriv0.mem", size12_type1_frame0_deriv0);
$readmemb("size12_type1_frame0_deriv1.mem", size12_type1_frame0_deriv1);
$readmemb("size12_type1_frame0_deriv2.mem", size12_type1_frame0_deriv2);
$readmemb("size12_type1_frame0_deriv3.mem", size12_type1_frame0_deriv3);
$readmemb("size12_type1_frame1_deriv0.mem", size12_type1_frame1_deriv0);
$readmemb("size12_type1_frame1_deriv1.mem", size12_type1_frame1_deriv1);
$readmemb("size12_type1_frame1_deriv2.mem", size12_type1_frame1_deriv2);
$readmemb("size12_type1_frame1_deriv3.mem", size12_type1_frame1_deriv3);
$readmemb("size13_type0_frame0_deriv0.mem", size13_type0_frame0_deriv0);
$readmemb("size13_type0_frame0_deriv1.mem", size13_type0_frame0_deriv1);
$readmemb("size13_type0_frame0_deriv2.mem", size13_type0_frame0_deriv2);
$readmemb("size13_type0_frame0_deriv3.mem", size13_type0_frame0_deriv3);
$readmemb("size13_type0_frame1_deriv0.mem", size13_type0_frame1_deriv0);
$readmemb("size13_type0_frame1_deriv1.mem", size13_type0_frame1_deriv1);
$readmemb("size13_type0_frame1_deriv2.mem", size13_type0_frame1_deriv2);
$readmemb("size13_type0_frame1_deriv3.mem", size13_type0_frame1_deriv3);
$readmemb("size13_type1_frame0_deriv0.mem", size13_type1_frame0_deriv0);
$readmemb("size13_type1_frame0_deriv1.mem", size13_type1_frame0_deriv1);
$readmemb("size13_type1_frame0_deriv2.mem", size13_type1_frame0_deriv2);
$readmemb("size13_type1_frame0_deriv3.mem", size13_type1_frame0_deriv3);
$readmemb("size13_type1_frame1_deriv0.mem", size13_type1_frame1_deriv0);
$readmemb("size13_type1_frame1_deriv1.mem", size13_type1_frame1_deriv1);
$readmemb("size13_type1_frame1_deriv2.mem", size13_type1_frame1_deriv2);
$readmemb("size13_type1_frame1_deriv3.mem", size13_type1_frame1_deriv3);
$readmemb("size14_type0_frame0_deriv0.mem", size14_type0_frame0_deriv0);
$readmemb("size14_type0_frame0_deriv1.mem", size14_type0_frame0_deriv1);
$readmemb("size14_type0_frame0_deriv2.mem", size14_type0_frame0_deriv2);
$readmemb("size14_type0_frame0_deriv3.mem", size14_type0_frame0_deriv3);
$readmemb("size14_type0_frame1_deriv0.mem", size14_type0_frame1_deriv0);
$readmemb("size14_type0_frame1_deriv1.mem", size14_type0_frame1_deriv1);
$readmemb("size14_type0_frame1_deriv2.mem", size14_type0_frame1_deriv2);
$readmemb("size14_type0_frame1_deriv3.mem", size14_type0_frame1_deriv3);
$readmemb("size14_type1_frame0_deriv0.mem", size14_type1_frame0_deriv0);
$readmemb("size14_type1_frame0_deriv1.mem", size14_type1_frame0_deriv1);
$readmemb("size14_type1_frame0_deriv2.mem", size14_type1_frame0_deriv2);
$readmemb("size14_type1_frame0_deriv3.mem", size14_type1_frame0_deriv3);
$readmemb("size14_type1_frame1_deriv0.mem", size14_type1_frame1_deriv0);
$readmemb("size14_type1_frame1_deriv1.mem", size14_type1_frame1_deriv1);
$readmemb("size14_type1_frame1_deriv2.mem", size14_type1_frame1_deriv2);
$readmemb("size14_type1_frame1_deriv3.mem", size14_type1_frame1_deriv3);
$readmemb("size15_type0_frame0_deriv0.mem", size15_type0_frame0_deriv0);
$readmemb("size15_type0_frame0_deriv1.mem", size15_type0_frame0_deriv1);
$readmemb("size15_type0_frame0_deriv2.mem", size15_type0_frame0_deriv2);
$readmemb("size15_type0_frame0_deriv3.mem", size15_type0_frame0_deriv3);
$readmemb("size15_type0_frame1_deriv0.mem", size15_type0_frame1_deriv0);
$readmemb("size15_type0_frame1_deriv1.mem", size15_type0_frame1_deriv1);
$readmemb("size15_type0_frame1_deriv2.mem", size15_type0_frame1_deriv2);
$readmemb("size15_type0_frame1_deriv3.mem", size15_type0_frame1_deriv3);
$readmemb("size15_type1_frame0_deriv0.mem", size15_type1_frame0_deriv0);
$readmemb("size15_type1_frame0_deriv1.mem", size15_type1_frame0_deriv1);
$readmemb("size15_type1_frame0_deriv2.mem", size15_type1_frame0_deriv2);
$readmemb("size15_type1_frame0_deriv3.mem", size15_type1_frame0_deriv3);
$readmemb("size15_type1_frame1_deriv0.mem", size15_type1_frame1_deriv0);
$readmemb("size15_type1_frame1_deriv1.mem", size15_type1_frame1_deriv1);
$readmemb("size15_type1_frame1_deriv2.mem", size15_type1_frame1_deriv2);
$readmemb("size15_type1_frame1_deriv3.mem", size15_type1_frame1_deriv3);
end

always @* begin
case({size_select, alien_type, frame_num, deriv_select})
10'b0000000000: palette_out = size0_type0_frame0_deriv0[pixel_addr];
10'b0000000001: palette_out = size0_type0_frame0_deriv1[pixel_addr];
10'b0000000010: palette_out = size0_type0_frame0_deriv2[pixel_addr];
10'b0000000011: palette_out = size0_type0_frame0_deriv3[pixel_addr];
10'b0000000100: palette_out = size0_type0_frame1_deriv0[pixel_addr];
10'b0000000101: palette_out = size0_type0_frame1_deriv1[pixel_addr];
10'b0000000110: palette_out = size0_type0_frame1_deriv2[pixel_addr];
10'b0000000111: palette_out = size0_type0_frame1_deriv3[pixel_addr];
10'b0000010000: palette_out = size0_type1_frame0_deriv0[pixel_addr];
10'b0000010001: palette_out = size0_type1_frame0_deriv1[pixel_addr];
10'b0000010010: palette_out = size0_type1_frame0_deriv2[pixel_addr];
10'b0000010011: palette_out = size0_type1_frame0_deriv3[pixel_addr];
10'b0000010100: palette_out = size0_type1_frame1_deriv0[pixel_addr];
10'b0000010101: palette_out = size0_type1_frame1_deriv1[pixel_addr];
10'b0000010110: palette_out = size0_type1_frame1_deriv2[pixel_addr];
10'b0000010111: palette_out = size0_type1_frame1_deriv3[pixel_addr];
10'b0001000000: palette_out = size1_type0_frame0_deriv0[pixel_addr];
10'b0001000001: palette_out = size1_type0_frame0_deriv1[pixel_addr];
10'b0001000010: palette_out = size1_type0_frame0_deriv2[pixel_addr];
10'b0001000011: palette_out = size1_type0_frame0_deriv3[pixel_addr];
10'b0001000100: palette_out = size1_type0_frame1_deriv0[pixel_addr];
10'b0001000101: palette_out = size1_type0_frame1_deriv1[pixel_addr];
10'b0001000110: palette_out = size1_type0_frame1_deriv2[pixel_addr];
10'b0001000111: palette_out = size1_type0_frame1_deriv3[pixel_addr];
10'b0001010000: palette_out = size1_type1_frame0_deriv0[pixel_addr];
10'b0001010001: palette_out = size1_type1_frame0_deriv1[pixel_addr];
10'b0001010010: palette_out = size1_type1_frame0_deriv2[pixel_addr];
10'b0001010011: palette_out = size1_type1_frame0_deriv3[pixel_addr];
10'b0001010100: palette_out = size1_type1_frame1_deriv0[pixel_addr];
10'b0001010101: palette_out = size1_type1_frame1_deriv1[pixel_addr];
10'b0001010110: palette_out = size1_type1_frame1_deriv2[pixel_addr];
10'b0001010111: palette_out = size1_type1_frame1_deriv3[pixel_addr];
10'b0010000000: palette_out = size2_type0_frame0_deriv0[pixel_addr];
10'b0010000001: palette_out = size2_type0_frame0_deriv1[pixel_addr];
10'b0010000010: palette_out = size2_type0_frame0_deriv2[pixel_addr];
10'b0010000011: palette_out = size2_type0_frame0_deriv3[pixel_addr];
10'b0010000100: palette_out = size2_type0_frame1_deriv0[pixel_addr];
10'b0010000101: palette_out = size2_type0_frame1_deriv1[pixel_addr];
10'b0010000110: palette_out = size2_type0_frame1_deriv2[pixel_addr];
10'b0010000111: palette_out = size2_type0_frame1_deriv3[pixel_addr];
10'b0010010000: palette_out = size2_type1_frame0_deriv0[pixel_addr];
10'b0010010001: palette_out = size2_type1_frame0_deriv1[pixel_addr];
10'b0010010010: palette_out = size2_type1_frame0_deriv2[pixel_addr];
10'b0010010011: palette_out = size2_type1_frame0_deriv3[pixel_addr];
10'b0010010100: palette_out = size2_type1_frame1_deriv0[pixel_addr];
10'b0010010101: palette_out = size2_type1_frame1_deriv1[pixel_addr];
10'b0010010110: palette_out = size2_type1_frame1_deriv2[pixel_addr];
10'b0010010111: palette_out = size2_type1_frame1_deriv3[pixel_addr];
10'b0011000000: palette_out = size3_type0_frame0_deriv0[pixel_addr];
10'b0011000001: palette_out = size3_type0_frame0_deriv1[pixel_addr];
10'b0011000010: palette_out = size3_type0_frame0_deriv2[pixel_addr];
10'b0011000011: palette_out = size3_type0_frame0_deriv3[pixel_addr];
10'b0011000100: palette_out = size3_type0_frame1_deriv0[pixel_addr];
10'b0011000101: palette_out = size3_type0_frame1_deriv1[pixel_addr];
10'b0011000110: palette_out = size3_type0_frame1_deriv2[pixel_addr];
10'b0011000111: palette_out = size3_type0_frame1_deriv3[pixel_addr];
10'b0011010000: palette_out = size3_type1_frame0_deriv0[pixel_addr];
10'b0011010001: palette_out = size3_type1_frame0_deriv1[pixel_addr];
10'b0011010010: palette_out = size3_type1_frame0_deriv2[pixel_addr];
10'b0011010011: palette_out = size3_type1_frame0_deriv3[pixel_addr];
10'b0011010100: palette_out = size3_type1_frame1_deriv0[pixel_addr];
10'b0011010101: palette_out = size3_type1_frame1_deriv1[pixel_addr];
10'b0011010110: palette_out = size3_type1_frame1_deriv2[pixel_addr];
10'b0011010111: palette_out = size3_type1_frame1_deriv3[pixel_addr];
10'b0100000000: palette_out = size4_type0_frame0_deriv0[pixel_addr];
10'b0100000001: palette_out = size4_type0_frame0_deriv1[pixel_addr];
10'b0100000010: palette_out = size4_type0_frame0_deriv2[pixel_addr];
10'b0100000011: palette_out = size4_type0_frame0_deriv3[pixel_addr];
10'b0100000100: palette_out = size4_type0_frame1_deriv0[pixel_addr];
10'b0100000101: palette_out = size4_type0_frame1_deriv1[pixel_addr];
10'b0100000110: palette_out = size4_type0_frame1_deriv2[pixel_addr];
10'b0100000111: palette_out = size4_type0_frame1_deriv3[pixel_addr];
10'b0100010000: palette_out = size4_type1_frame0_deriv0[pixel_addr];
10'b0100010001: palette_out = size4_type1_frame0_deriv1[pixel_addr];
10'b0100010010: palette_out = size4_type1_frame0_deriv2[pixel_addr];
10'b0100010011: palette_out = size4_type1_frame0_deriv3[pixel_addr];
10'b0100010100: palette_out = size4_type1_frame1_deriv0[pixel_addr];
10'b0100010101: palette_out = size4_type1_frame1_deriv1[pixel_addr];
10'b0100010110: palette_out = size4_type1_frame1_deriv2[pixel_addr];
10'b0100010111: palette_out = size4_type1_frame1_deriv3[pixel_addr];
10'b0101000000: palette_out = size5_type0_frame0_deriv0[pixel_addr];
10'b0101000001: palette_out = size5_type0_frame0_deriv1[pixel_addr];
10'b0101000010: palette_out = size5_type0_frame0_deriv2[pixel_addr];
10'b0101000011: palette_out = size5_type0_frame0_deriv3[pixel_addr];
10'b0101000100: palette_out = size5_type0_frame1_deriv0[pixel_addr];
10'b0101000101: palette_out = size5_type0_frame1_deriv1[pixel_addr];
10'b0101000110: palette_out = size5_type0_frame1_deriv2[pixel_addr];
10'b0101000111: palette_out = size5_type0_frame1_deriv3[pixel_addr];
10'b0101010000: palette_out = size5_type1_frame0_deriv0[pixel_addr];
10'b0101010001: palette_out = size5_type1_frame0_deriv1[pixel_addr];
10'b0101010010: palette_out = size5_type1_frame0_deriv2[pixel_addr];
10'b0101010011: palette_out = size5_type1_frame0_deriv3[pixel_addr];
10'b0101010100: palette_out = size5_type1_frame1_deriv0[pixel_addr];
10'b0101010101: palette_out = size5_type1_frame1_deriv1[pixel_addr];
10'b0101010110: palette_out = size5_type1_frame1_deriv2[pixel_addr];
10'b0101010111: palette_out = size5_type1_frame1_deriv3[pixel_addr];
10'b0110000000: palette_out = size6_type0_frame0_deriv0[pixel_addr];
10'b0110000001: palette_out = size6_type0_frame0_deriv1[pixel_addr];
10'b0110000010: palette_out = size6_type0_frame0_deriv2[pixel_addr];
10'b0110000011: palette_out = size6_type0_frame0_deriv3[pixel_addr];
10'b0110000100: palette_out = size6_type0_frame1_deriv0[pixel_addr];
10'b0110000101: palette_out = size6_type0_frame1_deriv1[pixel_addr];
10'b0110000110: palette_out = size6_type0_frame1_deriv2[pixel_addr];
10'b0110000111: palette_out = size6_type0_frame1_deriv3[pixel_addr];
10'b0110010000: palette_out = size6_type1_frame0_deriv0[pixel_addr];
10'b0110010001: palette_out = size6_type1_frame0_deriv1[pixel_addr];
10'b0110010010: palette_out = size6_type1_frame0_deriv2[pixel_addr];
10'b0110010011: palette_out = size6_type1_frame0_deriv3[pixel_addr];
10'b0110010100: palette_out = size6_type1_frame1_deriv0[pixel_addr];
10'b0110010101: palette_out = size6_type1_frame1_deriv1[pixel_addr];
10'b0110010110: palette_out = size6_type1_frame1_deriv2[pixel_addr];
10'b0110010111: palette_out = size6_type1_frame1_deriv3[pixel_addr];
10'b0111000000: palette_out = size7_type0_frame0_deriv0[pixel_addr];
10'b0111000001: palette_out = size7_type0_frame0_deriv1[pixel_addr];
10'b0111000010: palette_out = size7_type0_frame0_deriv2[pixel_addr];
10'b0111000011: palette_out = size7_type0_frame0_deriv3[pixel_addr];
10'b0111000100: palette_out = size7_type0_frame1_deriv0[pixel_addr];
10'b0111000101: palette_out = size7_type0_frame1_deriv1[pixel_addr];
10'b0111000110: palette_out = size7_type0_frame1_deriv2[pixel_addr];
10'b0111000111: palette_out = size7_type0_frame1_deriv3[pixel_addr];
10'b0111010000: palette_out = size7_type1_frame0_deriv0[pixel_addr];
10'b0111010001: palette_out = size7_type1_frame0_deriv1[pixel_addr];
10'b0111010010: palette_out = size7_type1_frame0_deriv2[pixel_addr];
10'b0111010011: palette_out = size7_type1_frame0_deriv3[pixel_addr];
10'b0111010100: palette_out = size7_type1_frame1_deriv0[pixel_addr];
10'b0111010101: palette_out = size7_type1_frame1_deriv1[pixel_addr];
10'b0111010110: palette_out = size7_type1_frame1_deriv2[pixel_addr];
10'b0111010111: palette_out = size7_type1_frame1_deriv3[pixel_addr];
10'b1000000000: palette_out = size8_type0_frame0_deriv0[pixel_addr];
10'b1000000001: palette_out = size8_type0_frame0_deriv1[pixel_addr];
10'b1000000010: palette_out = size8_type0_frame0_deriv2[pixel_addr];
10'b1000000011: palette_out = size8_type0_frame0_deriv3[pixel_addr];
10'b1000000100: palette_out = size8_type0_frame1_deriv0[pixel_addr];
10'b1000000101: palette_out = size8_type0_frame1_deriv1[pixel_addr];
10'b1000000110: palette_out = size8_type0_frame1_deriv2[pixel_addr];
10'b1000000111: palette_out = size8_type0_frame1_deriv3[pixel_addr];
10'b1000010000: palette_out = size8_type1_frame0_deriv0[pixel_addr];
10'b1000010001: palette_out = size8_type1_frame0_deriv1[pixel_addr];
10'b1000010010: palette_out = size8_type1_frame0_deriv2[pixel_addr];
10'b1000010011: palette_out = size8_type1_frame0_deriv3[pixel_addr];
10'b1000010100: palette_out = size8_type1_frame1_deriv0[pixel_addr];
10'b1000010101: palette_out = size8_type1_frame1_deriv1[pixel_addr];
10'b1000010110: palette_out = size8_type1_frame1_deriv2[pixel_addr];
10'b1000010111: palette_out = size8_type1_frame1_deriv3[pixel_addr];
10'b1001000000: palette_out = size9_type0_frame0_deriv0[pixel_addr];
10'b1001000001: palette_out = size9_type0_frame0_deriv1[pixel_addr];
10'b1001000010: palette_out = size9_type0_frame0_deriv2[pixel_addr];
10'b1001000011: palette_out = size9_type0_frame0_deriv3[pixel_addr];
10'b1001000100: palette_out = size9_type0_frame1_deriv0[pixel_addr];
10'b1001000101: palette_out = size9_type0_frame1_deriv1[pixel_addr];
10'b1001000110: palette_out = size9_type0_frame1_deriv2[pixel_addr];
10'b1001000111: palette_out = size9_type0_frame1_deriv3[pixel_addr];
10'b1001010000: palette_out = size9_type1_frame0_deriv0[pixel_addr];
10'b1001010001: palette_out = size9_type1_frame0_deriv1[pixel_addr];
10'b1001010010: palette_out = size9_type1_frame0_deriv2[pixel_addr];
10'b1001010011: palette_out = size9_type1_frame0_deriv3[pixel_addr];
10'b1001010100: palette_out = size9_type1_frame1_deriv0[pixel_addr];
10'b1001010101: palette_out = size9_type1_frame1_deriv1[pixel_addr];
10'b1001010110: palette_out = size9_type1_frame1_deriv2[pixel_addr];
10'b1001010111: palette_out = size9_type1_frame1_deriv3[pixel_addr];
10'b1010000000: palette_out = size10_type0_frame0_deriv0[pixel_addr];
10'b1010000001: palette_out = size10_type0_frame0_deriv1[pixel_addr];
10'b1010000010: palette_out = size10_type0_frame0_deriv2[pixel_addr];
10'b1010000011: palette_out = size10_type0_frame0_deriv3[pixel_addr];
10'b1010000100: palette_out = size10_type0_frame1_deriv0[pixel_addr];
10'b1010000101: palette_out = size10_type0_frame1_deriv1[pixel_addr];
10'b1010000110: palette_out = size10_type0_frame1_deriv2[pixel_addr];
10'b1010000111: palette_out = size10_type0_frame1_deriv3[pixel_addr];
10'b1010010000: palette_out = size10_type1_frame0_deriv0[pixel_addr];
10'b1010010001: palette_out = size10_type1_frame0_deriv1[pixel_addr];
10'b1010010010: palette_out = size10_type1_frame0_deriv2[pixel_addr];
10'b1010010011: palette_out = size10_type1_frame0_deriv3[pixel_addr];
10'b1010010100: palette_out = size10_type1_frame1_deriv0[pixel_addr];
10'b1010010101: palette_out = size10_type1_frame1_deriv1[pixel_addr];
10'b1010010110: palette_out = size10_type1_frame1_deriv2[pixel_addr];
10'b1010010111: palette_out = size10_type1_frame1_deriv3[pixel_addr];
10'b1011000000: palette_out = size11_type0_frame0_deriv0[pixel_addr];
10'b1011000001: palette_out = size11_type0_frame0_deriv1[pixel_addr];
10'b1011000010: palette_out = size11_type0_frame0_deriv2[pixel_addr];
10'b1011000011: palette_out = size11_type0_frame0_deriv3[pixel_addr];
10'b1011000100: palette_out = size11_type0_frame1_deriv0[pixel_addr];
10'b1011000101: palette_out = size11_type0_frame1_deriv1[pixel_addr];
10'b1011000110: palette_out = size11_type0_frame1_deriv2[pixel_addr];
10'b1011000111: palette_out = size11_type0_frame1_deriv3[pixel_addr];
10'b1011010000: palette_out = size11_type1_frame0_deriv0[pixel_addr];
10'b1011010001: palette_out = size11_type1_frame0_deriv1[pixel_addr];
10'b1011010010: palette_out = size11_type1_frame0_deriv2[pixel_addr];
10'b1011010011: palette_out = size11_type1_frame0_deriv3[pixel_addr];
10'b1011010100: palette_out = size11_type1_frame1_deriv0[pixel_addr];
10'b1011010101: palette_out = size11_type1_frame1_deriv1[pixel_addr];
10'b1011010110: palette_out = size11_type1_frame1_deriv2[pixel_addr];
10'b1011010111: palette_out = size11_type1_frame1_deriv3[pixel_addr];
10'b1100000000: palette_out = size12_type0_frame0_deriv0[pixel_addr];
10'b1100000001: palette_out = size12_type0_frame0_deriv1[pixel_addr];
10'b1100000010: palette_out = size12_type0_frame0_deriv2[pixel_addr];
10'b1100000011: palette_out = size12_type0_frame0_deriv3[pixel_addr];
10'b1100000100: palette_out = size12_type0_frame1_deriv0[pixel_addr];
10'b1100000101: palette_out = size12_type0_frame1_deriv1[pixel_addr];
10'b1100000110: palette_out = size12_type0_frame1_deriv2[pixel_addr];
10'b1100000111: palette_out = size12_type0_frame1_deriv3[pixel_addr];
10'b1100010000: palette_out = size12_type1_frame0_deriv0[pixel_addr];
10'b1100010001: palette_out = size12_type1_frame0_deriv1[pixel_addr];
10'b1100010010: palette_out = size12_type1_frame0_deriv2[pixel_addr];
10'b1100010011: palette_out = size12_type1_frame0_deriv3[pixel_addr];
10'b1100010100: palette_out = size12_type1_frame1_deriv0[pixel_addr];
10'b1100010101: palette_out = size12_type1_frame1_deriv1[pixel_addr];
10'b1100010110: palette_out = size12_type1_frame1_deriv2[pixel_addr];
10'b1100010111: palette_out = size12_type1_frame1_deriv3[pixel_addr];
10'b1101000000: palette_out = size13_type0_frame0_deriv0[pixel_addr];
10'b1101000001: palette_out = size13_type0_frame0_deriv1[pixel_addr];
10'b1101000010: palette_out = size13_type0_frame0_deriv2[pixel_addr];
10'b1101000011: palette_out = size13_type0_frame0_deriv3[pixel_addr];
10'b1101000100: palette_out = size13_type0_frame1_deriv0[pixel_addr];
10'b1101000101: palette_out = size13_type0_frame1_deriv1[pixel_addr];
10'b1101000110: palette_out = size13_type0_frame1_deriv2[pixel_addr];
10'b1101000111: palette_out = size13_type0_frame1_deriv3[pixel_addr];
10'b1101010000: palette_out = size13_type1_frame0_deriv0[pixel_addr];
10'b1101010001: palette_out = size13_type1_frame0_deriv1[pixel_addr];
10'b1101010010: palette_out = size13_type1_frame0_deriv2[pixel_addr];
10'b1101010011: palette_out = size13_type1_frame0_deriv3[pixel_addr];
10'b1101010100: palette_out = size13_type1_frame1_deriv0[pixel_addr];
10'b1101010101: palette_out = size13_type1_frame1_deriv1[pixel_addr];
10'b1101010110: palette_out = size13_type1_frame1_deriv2[pixel_addr];
10'b1101010111: palette_out = size13_type1_frame1_deriv3[pixel_addr];
10'b1110000000: palette_out = size14_type0_frame0_deriv0[pixel_addr];
10'b1110000001: palette_out = size14_type0_frame0_deriv1[pixel_addr];
10'b1110000010: palette_out = size14_type0_frame0_deriv2[pixel_addr];
10'b1110000011: palette_out = size14_type0_frame0_deriv3[pixel_addr];
10'b1110000100: palette_out = size14_type0_frame1_deriv0[pixel_addr];
10'b1110000101: palette_out = size14_type0_frame1_deriv1[pixel_addr];
10'b1110000110: palette_out = size14_type0_frame1_deriv2[pixel_addr];
10'b1110000111: palette_out = size14_type0_frame1_deriv3[pixel_addr];
10'b1110010000: palette_out = size14_type1_frame0_deriv0[pixel_addr];
10'b1110010001: palette_out = size14_type1_frame0_deriv1[pixel_addr];
10'b1110010010: palette_out = size14_type1_frame0_deriv2[pixel_addr];
10'b1110010011: palette_out = size14_type1_frame0_deriv3[pixel_addr];
10'b1110010100: palette_out = size14_type1_frame1_deriv0[pixel_addr];
10'b1110010101: palette_out = size14_type1_frame1_deriv1[pixel_addr];
10'b1110010110: palette_out = size14_type1_frame1_deriv2[pixel_addr];
10'b1110010111: palette_out = size14_type1_frame1_deriv3[pixel_addr];
10'b1111000000: palette_out = size15_type0_frame0_deriv0[pixel_addr];
10'b1111000001: palette_out = size15_type0_frame0_deriv1[pixel_addr];
10'b1111000010: palette_out = size15_type0_frame0_deriv2[pixel_addr];
10'b1111000011: palette_out = size15_type0_frame0_deriv3[pixel_addr];
10'b1111000100: palette_out = size15_type0_frame1_deriv0[pixel_addr];
10'b1111000101: palette_out = size15_type0_frame1_deriv1[pixel_addr];
10'b1111000110: palette_out = size15_type0_frame1_deriv2[pixel_addr];
10'b1111000111: palette_out = size15_type0_frame1_deriv3[pixel_addr];
10'b1111010000: palette_out = size15_type1_frame0_deriv0[pixel_addr];
10'b1111010001: palette_out = size15_type1_frame0_deriv1[pixel_addr];
10'b1111010010: palette_out = size15_type1_frame0_deriv2[pixel_addr];
10'b1111010011: palette_out = size15_type1_frame0_deriv3[pixel_addr];
10'b1111010100: palette_out = size15_type1_frame1_deriv0[pixel_addr];
10'b1111010101: palette_out = size15_type1_frame1_deriv1[pixel_addr];
10'b1111010110: palette_out = size15_type1_frame1_deriv2[pixel_addr];
10'b1111010111: palette_out = size15_type1_frame1_deriv3[pixel_addr];
default : palette_out = 0;
endcase
end
    
endmodule
